magic
tech sky130A
magscale 1 2
timestamp 1756673146
<< viali >>
rect 121 3009 155 3043
rect 2973 3009 3007 3043
rect 397 2941 431 2975
rect 857 2941 891 2975
rect 1133 2941 1167 2975
rect 2605 2941 2639 2975
rect 2789 2941 2823 2975
rect 3157 2805 3191 2839
rect 397 2465 431 2499
rect 857 2465 891 2499
rect 1133 2465 1167 2499
rect 2605 2465 2639 2499
rect 2789 2465 2823 2499
rect 121 2397 155 2431
rect 2973 2397 3007 2431
rect 3157 2261 3191 2295
rect 121 1921 155 1955
rect 2973 1921 3007 1955
rect 397 1853 431 1887
rect 857 1853 891 1887
rect 1133 1853 1167 1887
rect 2605 1853 2639 1887
rect 2789 1853 2823 1887
rect 3157 1717 3191 1751
rect 857 1377 891 1411
rect 1133 1377 1167 1411
rect 2605 1377 2639 1411
rect 2789 1377 2823 1411
rect 2973 1309 3007 1343
rect 3157 1173 3191 1207
rect 2973 833 3007 867
rect 857 765 891 799
rect 1133 765 1167 799
rect 2605 765 2639 799
rect 2789 765 2823 799
rect 3157 629 3191 663
rect 673 357 707 391
rect 857 289 891 323
rect 1133 289 1167 323
rect 2605 289 2639 323
rect 2789 289 2823 323
rect 29 221 63 255
rect 2973 221 3007 255
rect 3157 85 3191 119
<< metal1 >>
rect 750 3068 756 3120
rect 808 3108 814 3120
rect 808 3080 1624 3108
rect 808 3068 814 3080
rect 106 3000 112 3052
rect 164 3000 170 3052
rect 2958 3000 2964 3052
rect 3016 3000 3022 3052
rect 385 2975 443 2981
rect 385 2941 397 2975
rect 431 2972 443 2975
rect 842 2972 848 2984
rect 431 2944 848 2972
rect 431 2941 443 2944
rect 385 2935 443 2941
rect 842 2932 848 2944
rect 900 2932 906 2984
rect 1121 2975 1179 2981
rect 1121 2941 1133 2975
rect 1167 2972 1179 2975
rect 1854 2972 1860 2984
rect 1167 2944 1860 2972
rect 1167 2941 1179 2944
rect 1121 2935 1179 2941
rect 1854 2932 1860 2944
rect 1912 2932 1918 2984
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2639 2944 2789 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 2777 2941 2789 2944
rect 2823 2972 2835 2975
rect 3510 2972 3516 2984
rect 2823 2944 3516 2972
rect 2823 2941 2835 2944
rect 2777 2935 2835 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3142 2796 3148 2848
rect 3200 2796 3206 2848
rect 385 2499 443 2505
rect 385 2465 397 2499
rect 431 2496 443 2499
rect 750 2496 756 2508
rect 431 2468 756 2496
rect 431 2465 443 2468
rect 385 2459 443 2465
rect 750 2456 756 2468
rect 808 2456 814 2508
rect 842 2456 848 2508
rect 900 2456 906 2508
rect 1121 2499 1179 2505
rect 1121 2465 1133 2499
rect 1167 2496 1179 2499
rect 1762 2496 1768 2508
rect 1167 2468 1768 2496
rect 1167 2465 1179 2468
rect 1121 2459 1179 2465
rect 1762 2456 1768 2468
rect 1820 2456 1826 2508
rect 1854 2456 1860 2508
rect 1912 2496 1918 2508
rect 2593 2499 2651 2505
rect 2593 2496 2605 2499
rect 1912 2468 2605 2496
rect 1912 2456 1918 2468
rect 2593 2465 2605 2468
rect 2639 2496 2651 2499
rect 2777 2499 2835 2505
rect 2777 2496 2789 2499
rect 2639 2468 2789 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 2777 2465 2789 2468
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 106 2388 112 2440
rect 164 2388 170 2440
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 750 2320 756 2372
rect 808 2360 814 2372
rect 808 2332 1624 2360
rect 808 2320 814 2332
rect 3142 2252 3148 2304
rect 3200 2252 3206 2304
rect 2958 2088 2964 2100
rect 400 2060 2964 2088
rect 106 1912 112 1964
rect 164 1912 170 1964
rect 400 1899 428 2060
rect 2958 2048 2964 2060
rect 3016 2048 3022 2100
rect 750 1980 756 2032
rect 808 2020 814 2032
rect 808 1992 1624 2020
rect 808 1980 814 1992
rect 2958 1912 2964 1964
rect 3016 1912 3022 1964
rect 391 1887 437 1899
rect 391 1853 397 1887
rect 431 1853 437 1887
rect 391 1841 437 1853
rect 842 1844 848 1896
rect 900 1844 906 1896
rect 1121 1887 1179 1893
rect 1121 1853 1133 1887
rect 1167 1884 1179 1887
rect 1670 1884 1676 1896
rect 1167 1856 1676 1884
rect 1167 1853 1179 1856
rect 1121 1847 1179 1853
rect 1670 1844 1676 1856
rect 1728 1844 1734 1896
rect 1762 1844 1768 1896
rect 1820 1884 1826 1896
rect 2593 1887 2651 1893
rect 2593 1884 2605 1887
rect 1820 1856 2605 1884
rect 1820 1844 1826 1856
rect 2593 1853 2605 1856
rect 2639 1884 2651 1887
rect 2777 1887 2835 1893
rect 2777 1884 2789 1887
rect 2639 1856 2789 1884
rect 2639 1853 2651 1856
rect 2593 1847 2651 1853
rect 2777 1853 2789 1856
rect 2823 1853 2835 1887
rect 2777 1847 2835 1853
rect 3142 1708 3148 1760
rect 3200 1708 3206 1760
rect 842 1368 848 1420
rect 900 1368 906 1420
rect 1121 1411 1179 1417
rect 1121 1377 1133 1411
rect 1167 1408 1179 1411
rect 1578 1408 1584 1420
rect 1167 1380 1584 1408
rect 1167 1377 1179 1380
rect 1121 1371 1179 1377
rect 1578 1368 1584 1380
rect 1636 1368 1642 1420
rect 1670 1368 1676 1420
rect 1728 1408 1734 1420
rect 2593 1411 2651 1417
rect 2593 1408 2605 1411
rect 1728 1380 2605 1408
rect 1728 1368 1734 1380
rect 2593 1377 2605 1380
rect 2639 1408 2651 1411
rect 2777 1411 2835 1417
rect 2777 1408 2789 1411
rect 2639 1380 2789 1408
rect 2639 1377 2651 1380
rect 2593 1371 2651 1377
rect 2777 1377 2789 1380
rect 2823 1377 2835 1411
rect 2777 1371 2835 1377
rect 2958 1300 2964 1352
rect 3016 1300 3022 1352
rect 750 1232 756 1284
rect 808 1272 814 1284
rect 808 1244 1624 1272
rect 808 1232 814 1244
rect 3142 1164 3148 1216
rect 3200 1164 3206 1216
rect 750 892 756 944
rect 808 932 814 944
rect 808 904 1624 932
rect 808 892 814 904
rect 2958 824 2964 876
rect 3016 824 3022 876
rect 842 756 848 808
rect 900 756 906 808
rect 1121 799 1179 805
rect 1121 765 1133 799
rect 1167 796 1179 799
rect 1486 796 1492 808
rect 1167 768 1492 796
rect 1167 765 1179 768
rect 1121 759 1179 765
rect 1486 756 1492 768
rect 1544 756 1550 808
rect 1578 756 1584 808
rect 1636 796 1642 808
rect 2593 799 2651 805
rect 2593 796 2605 799
rect 1636 768 2605 796
rect 1636 756 1642 768
rect 2593 765 2605 768
rect 2639 796 2651 799
rect 2777 799 2835 805
rect 2777 796 2789 799
rect 2639 768 2789 796
rect 2639 765 2651 768
rect 2593 759 2651 765
rect 2777 765 2789 768
rect 2823 765 2835 799
rect 2777 759 2835 765
rect 3142 620 3148 672
rect 3200 620 3206 672
rect 661 391 719 397
rect 661 357 673 391
rect 707 388 719 391
rect 707 360 980 388
rect 707 357 719 360
rect 661 351 719 357
rect 842 280 848 332
rect 900 280 906 332
rect 952 320 980 360
rect 1121 323 1179 329
rect 1121 320 1133 323
rect 952 292 1133 320
rect 1121 289 1133 292
rect 1167 289 1179 323
rect 1121 283 1179 289
rect 1486 280 1492 332
rect 1544 320 1550 332
rect 2593 323 2651 329
rect 2593 320 2605 323
rect 1544 292 2605 320
rect 1544 280 1550 292
rect 2593 289 2605 292
rect 2639 320 2651 323
rect 2777 323 2835 329
rect 2777 320 2789 323
rect 2639 292 2789 320
rect 2639 289 2651 292
rect 2593 283 2651 289
rect 2777 289 2789 292
rect 2823 289 2835 323
rect 2777 283 2835 289
rect 13 255 79 261
rect 13 252 29 255
rect 0 224 29 252
rect 13 221 29 224
rect 63 221 79 255
rect 13 215 79 221
rect 2958 212 2964 264
rect 3016 212 3022 264
rect 3510 212 3516 264
rect 3568 252 3574 264
rect 3568 224 3680 252
rect 3568 212 3574 224
rect 750 144 756 196
rect 808 184 814 196
rect 808 156 1624 184
rect 808 144 814 156
rect 3142 76 3148 128
rect 3200 76 3206 128
<< via1 >>
rect 340 3222 580 3306
rect 756 3068 808 3120
rect 112 3043 164 3052
rect 112 3009 121 3043
rect 121 3009 155 3043
rect 155 3009 164 3043
rect 112 3000 164 3009
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 848 2975 900 2984
rect 848 2941 857 2975
rect 857 2941 891 2975
rect 891 2941 900 2975
rect 848 2932 900 2941
rect 1860 2932 1912 2984
rect 3516 2932 3568 2984
rect 3148 2839 3200 2848
rect 3148 2805 3157 2839
rect 3157 2805 3191 2839
rect 3191 2805 3200 2839
rect 3148 2796 3200 2805
rect 20 2678 260 2762
rect 756 2456 808 2508
rect 848 2499 900 2508
rect 848 2465 857 2499
rect 857 2465 891 2499
rect 891 2465 900 2499
rect 848 2456 900 2465
rect 1768 2456 1820 2508
rect 1860 2456 1912 2508
rect 112 2431 164 2440
rect 112 2397 121 2431
rect 121 2397 155 2431
rect 155 2397 164 2431
rect 112 2388 164 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 756 2320 808 2372
rect 3148 2295 3200 2304
rect 3148 2261 3157 2295
rect 3157 2261 3191 2295
rect 3191 2261 3200 2295
rect 3148 2252 3200 2261
rect 340 2134 580 2218
rect 112 1955 164 1964
rect 112 1921 121 1955
rect 121 1921 155 1955
rect 155 1921 164 1955
rect 112 1912 164 1921
rect 2964 2048 3016 2100
rect 756 1980 808 2032
rect 2964 1955 3016 1964
rect 2964 1921 2973 1955
rect 2973 1921 3007 1955
rect 3007 1921 3016 1955
rect 2964 1912 3016 1921
rect 848 1887 900 1896
rect 848 1853 857 1887
rect 857 1853 891 1887
rect 891 1853 900 1887
rect 848 1844 900 1853
rect 1676 1844 1728 1896
rect 1768 1844 1820 1896
rect 3148 1751 3200 1760
rect 3148 1717 3157 1751
rect 3157 1717 3191 1751
rect 3191 1717 3200 1751
rect 3148 1708 3200 1717
rect 20 1590 260 1674
rect 848 1411 900 1420
rect 848 1377 857 1411
rect 857 1377 891 1411
rect 891 1377 900 1411
rect 848 1368 900 1377
rect 1584 1368 1636 1420
rect 1676 1368 1728 1420
rect 2964 1343 3016 1352
rect 2964 1309 2973 1343
rect 2973 1309 3007 1343
rect 3007 1309 3016 1343
rect 2964 1300 3016 1309
rect 756 1232 808 1284
rect 3148 1207 3200 1216
rect 3148 1173 3157 1207
rect 3157 1173 3191 1207
rect 3191 1173 3200 1207
rect 3148 1164 3200 1173
rect 340 1046 580 1130
rect 756 892 808 944
rect 2964 867 3016 876
rect 2964 833 2973 867
rect 2973 833 3007 867
rect 3007 833 3016 867
rect 2964 824 3016 833
rect 848 799 900 808
rect 848 765 857 799
rect 857 765 891 799
rect 891 765 900 799
rect 848 756 900 765
rect 1492 756 1544 808
rect 1584 756 1636 808
rect 3148 663 3200 672
rect 3148 629 3157 663
rect 3157 629 3191 663
rect 3191 629 3200 663
rect 3148 620 3200 629
rect 20 502 260 586
rect 848 323 900 332
rect 848 289 857 323
rect 857 289 891 323
rect 891 289 900 323
rect 848 280 900 289
rect 1492 280 1544 332
rect 2964 255 3016 264
rect 2964 221 2973 255
rect 2973 221 3007 255
rect 3007 221 3016 255
rect 2964 212 3016 221
rect 3516 212 3568 264
rect 756 144 808 196
rect 3148 119 3200 128
rect 3148 85 3157 119
rect 3157 85 3191 119
rect 3191 85 3200 119
rect 3148 76 3200 85
rect 340 -42 580 42
<< metal2 >>
rect 340 3306 580 3312
rect 340 3216 580 3222
rect 756 3120 808 3126
rect 756 3062 808 3068
rect 110 3052 166 3058
rect 110 3020 112 3052
rect 164 3020 166 3052
rect 110 2955 166 2964
rect 20 2762 260 2768
rect 20 2672 260 2678
rect 768 2514 796 3062
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 848 2984 900 2990
rect 848 2926 900 2932
rect 1860 2984 1912 2990
rect 1860 2926 1912 2932
rect 860 2514 888 2926
rect 1872 2514 1900 2926
rect 756 2508 808 2514
rect 110 2476 166 2485
rect 756 2450 808 2456
rect 848 2508 900 2514
rect 848 2450 900 2456
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 110 2388 112 2420
rect 164 2388 166 2420
rect 110 2382 166 2388
rect 768 2378 796 2450
rect 756 2372 808 2378
rect 756 2314 808 2320
rect 340 2218 580 2224
rect 340 2128 580 2134
rect 768 2038 796 2314
rect 756 2032 808 2038
rect 756 1974 808 1980
rect 110 1964 166 1970
rect 110 1932 112 1964
rect 164 1932 166 1964
rect 110 1867 166 1876
rect 20 1674 260 1680
rect 20 1584 260 1590
rect 768 1290 796 1974
rect 860 1902 888 2450
rect 1780 1902 1808 2450
rect 2976 2446 3004 2994
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3146 2850 3202 2859
rect 3146 2785 3202 2794
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2976 2106 3004 2382
rect 3146 2306 3202 2315
rect 3146 2241 3202 2250
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 2976 1970 3004 2042
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 848 1896 900 1902
rect 848 1838 900 1844
rect 1676 1896 1728 1902
rect 1676 1838 1728 1844
rect 1768 1896 1820 1902
rect 1768 1838 1820 1844
rect 860 1426 888 1838
rect 1688 1426 1716 1838
rect 848 1420 900 1426
rect 848 1362 900 1368
rect 1584 1420 1636 1426
rect 1584 1362 1636 1368
rect 1676 1420 1728 1426
rect 1676 1362 1728 1368
rect 756 1284 808 1290
rect 756 1226 808 1232
rect 340 1130 580 1136
rect 340 1040 580 1046
rect 768 950 796 1226
rect 756 944 808 950
rect 756 886 808 892
rect 20 586 260 592
rect 20 496 260 502
rect 768 202 796 886
rect 860 814 888 1362
rect 1596 814 1624 1362
rect 2976 1358 3004 1906
rect 3146 1762 3202 1771
rect 3146 1697 3202 1706
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 2976 882 3004 1294
rect 3146 1218 3202 1227
rect 3146 1153 3202 1162
rect 2964 876 3016 882
rect 2964 818 3016 824
rect 848 808 900 814
rect 848 750 900 756
rect 1492 808 1544 814
rect 1492 750 1544 756
rect 1584 808 1636 814
rect 1584 750 1636 756
rect 860 338 888 750
rect 1504 338 1532 750
rect 848 332 900 338
rect 848 274 900 280
rect 1492 332 1544 338
rect 1492 274 1544 280
rect 2976 270 3004 818
rect 3146 674 3202 683
rect 3146 609 3202 618
rect 3528 270 3556 2926
rect 2964 264 3016 270
rect 2964 206 3016 212
rect 3516 264 3568 270
rect 3516 206 3568 212
rect 756 196 808 202
rect 756 138 808 144
rect 3146 130 3202 139
rect 3146 65 3202 74
rect 340 42 580 48
rect 340 -48 580 -42
<< via2 >>
rect 345 3225 575 3303
rect 110 3000 112 3020
rect 112 3000 164 3020
rect 164 3000 166 3020
rect 110 2964 166 3000
rect 25 2681 255 2759
rect 110 2440 166 2476
rect 110 2420 112 2440
rect 112 2420 164 2440
rect 164 2420 166 2440
rect 345 2137 575 2215
rect 110 1912 112 1932
rect 112 1912 164 1932
rect 164 1912 166 1932
rect 110 1876 166 1912
rect 25 1593 255 1671
rect 3146 2848 3202 2850
rect 3146 2796 3148 2848
rect 3148 2796 3200 2848
rect 3200 2796 3202 2848
rect 3146 2794 3202 2796
rect 3146 2304 3202 2306
rect 3146 2252 3148 2304
rect 3148 2252 3200 2304
rect 3200 2252 3202 2304
rect 3146 2250 3202 2252
rect 345 1049 575 1127
rect 25 505 255 583
rect 3146 1760 3202 1762
rect 3146 1708 3148 1760
rect 3148 1708 3200 1760
rect 3200 1708 3202 1760
rect 3146 1706 3202 1708
rect 3146 1216 3202 1218
rect 3146 1164 3148 1216
rect 3148 1164 3200 1216
rect 3200 1164 3202 1216
rect 3146 1162 3202 1164
rect 3146 672 3202 674
rect 3146 620 3148 672
rect 3148 620 3200 672
rect 3200 620 3202 672
rect 3146 618 3202 620
rect 3146 128 3202 130
rect 3146 76 3148 128
rect 3148 76 3200 128
rect 3200 76 3202 128
rect 3146 74 3202 76
rect 345 -39 575 39
<< metal3 >>
rect 340 3306 580 3312
rect 340 3222 341 3306
rect 579 3222 580 3306
rect 340 3216 580 3222
rect 105 3022 171 3025
rect 0 3020 3680 3022
rect 0 2964 110 3020
rect 166 2964 3680 3020
rect 0 2962 3680 2964
rect 105 2959 171 2962
rect 996 2790 1002 2854
rect 1066 2852 1072 2854
rect 3141 2852 3207 2855
rect 1066 2850 3207 2852
rect 1066 2794 3146 2850
rect 3202 2794 3207 2850
rect 1066 2792 3207 2794
rect 1066 2790 1072 2792
rect 3141 2789 3207 2792
rect 20 2762 260 2768
rect 20 2678 21 2762
rect 259 2678 260 2762
rect 20 2672 260 2678
rect 105 2478 171 2481
rect 0 2476 3680 2478
rect 0 2420 110 2476
rect 166 2420 3680 2476
rect 0 2418 3680 2420
rect 105 2415 171 2418
rect 1115 2246 1121 2310
rect 1185 2308 1191 2310
rect 3141 2308 3207 2311
rect 1185 2306 3207 2308
rect 1185 2250 3146 2306
rect 3202 2250 3207 2306
rect 1185 2248 3207 2250
rect 1185 2246 1191 2248
rect 3141 2245 3207 2248
rect 340 2218 580 2224
rect 340 2134 341 2218
rect 579 2134 580 2218
rect 340 2128 580 2134
rect 105 1934 171 1937
rect 0 1932 3680 1934
rect 0 1876 110 1932
rect 166 1876 3680 1932
rect 0 1874 3680 1876
rect 105 1871 171 1874
rect 1235 1702 1241 1766
rect 1305 1764 1311 1766
rect 3141 1764 3207 1767
rect 1305 1762 3207 1764
rect 1305 1706 3146 1762
rect 3202 1706 3207 1762
rect 1305 1704 3207 1706
rect 1305 1702 1311 1704
rect 3141 1701 3207 1704
rect 20 1674 260 1680
rect 20 1590 21 1674
rect 259 1590 260 1674
rect 20 1584 260 1590
rect 1355 1158 1361 1222
rect 1425 1220 1431 1222
rect 3141 1220 3207 1223
rect 1425 1218 3207 1220
rect 1425 1162 3146 1218
rect 3202 1162 3207 1218
rect 1425 1160 3207 1162
rect 1425 1158 1431 1160
rect 3141 1157 3207 1160
rect 340 1130 580 1136
rect 340 1046 341 1130
rect 579 1046 580 1130
rect 340 1040 580 1046
rect 1475 614 1481 678
rect 1545 676 1551 678
rect 3141 676 3207 679
rect 1545 674 3207 676
rect 1545 618 3146 674
rect 3202 618 3207 674
rect 1545 616 3207 618
rect 1545 614 1551 616
rect 3141 613 3207 616
rect 20 586 260 592
rect 20 502 21 586
rect 259 502 260 586
rect 20 496 260 502
rect 1595 70 1601 134
rect 1665 132 1671 134
rect 3141 132 3207 135
rect 1665 130 3207 132
rect 1665 74 3146 130
rect 3202 74 3207 130
rect 1665 72 3207 74
rect 1665 70 1671 72
rect 3141 69 3207 72
rect 340 42 580 48
rect 340 -42 341 42
rect 579 -42 580 42
rect 340 -48 580 -42
<< via3 >>
rect 341 3303 579 3306
rect 341 3225 345 3303
rect 345 3225 575 3303
rect 575 3225 579 3303
rect 341 3222 579 3225
rect 1002 2790 1066 2854
rect 21 2759 259 2762
rect 21 2681 25 2759
rect 25 2681 255 2759
rect 255 2681 259 2759
rect 21 2678 259 2681
rect 1121 2246 1185 2310
rect 341 2215 579 2218
rect 341 2137 345 2215
rect 345 2137 575 2215
rect 575 2137 579 2215
rect 341 2134 579 2137
rect 1241 1702 1305 1766
rect 21 1671 259 1674
rect 21 1593 25 1671
rect 25 1593 255 1671
rect 255 1593 259 1671
rect 21 1590 259 1593
rect 1361 1158 1425 1222
rect 341 1127 579 1130
rect 341 1049 345 1127
rect 345 1049 575 1127
rect 575 1049 579 1127
rect 341 1046 579 1049
rect 1481 614 1545 678
rect 21 583 259 586
rect 21 505 25 583
rect 25 505 255 583
rect 255 505 259 583
rect 21 502 259 505
rect 1601 70 1665 134
rect 341 39 579 42
rect 341 -39 345 39
rect 345 -39 575 39
rect 575 -39 579 39
rect 341 -42 579 -39
<< metal4 >>
rect 20 2762 260 3312
rect 20 2678 21 2762
rect 259 2678 260 2762
rect 20 1674 260 2678
rect 20 1590 21 1674
rect 259 1590 260 1674
rect 20 586 260 1590
rect 20 502 21 586
rect 259 502 260 586
rect 20 -48 260 502
rect 340 3306 580 3312
rect 340 3222 341 3306
rect 579 3222 580 3306
rect 340 2218 580 3222
rect 1001 2854 1067 2855
rect 1001 2834 1002 2854
rect 340 2134 341 2218
rect 579 2134 580 2218
rect 340 1130 580 2134
rect 340 1046 341 1130
rect 579 1046 580 1130
rect 340 42 580 1046
rect 340 -42 341 42
rect 579 -42 580 42
rect 340 -48 580 -42
rect 1000 2790 1002 2834
rect 1066 2790 1067 2854
rect 1000 2789 1067 2790
rect 1000 2781 1061 2789
rect 1000 -48 1060 2781
rect 1120 2310 1186 2311
rect 1120 2246 1121 2310
rect 1185 2246 1186 2310
rect 1120 2245 1186 2246
rect 1120 -48 1180 2245
rect 1240 1766 1306 1767
rect 1240 1702 1241 1766
rect 1305 1702 1306 1766
rect 1240 1701 1306 1702
rect 1240 -48 1300 1701
rect 1360 1222 1426 1223
rect 1360 1158 1361 1222
rect 1425 1158 1426 1222
rect 1360 1157 1426 1158
rect 1360 -48 1420 1157
rect 1480 678 1546 679
rect 1480 614 1481 678
rect 1545 614 1546 678
rect 1480 613 1546 614
rect 1480 -48 1540 613
rect 1600 134 1666 135
rect 1600 70 1601 134
rect 1665 70 1666 134
rect 1600 69 1666 70
rect 1600 -48 1660 69
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 2760 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_1
timestamp 1755005639
transform 1 0 2760 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_2
timestamp 1755005639
transform 1 0 2760 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_3
timestamp 1755005639
transform 1 0 2760 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_4
timestamp 1755005639
transform 1 0 2760 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_5
timestamp 1755005639
transform 1 0 2760 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 0 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_1
timestamp 1755005639
transform 1 0 0 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_2
timestamp 1755005639
transform 1 0 0 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s50_2  sky130_fd_sc_hd__clkdlybuf4s50_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 0 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 552 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1755005639
transform 1 0 552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1755005639
transform 1 0 552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 3312 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1755005639
transform 1 0 3312 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1755005639
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1755005639
transform 1 0 3312 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1755005639
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1755005639
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 0 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1755005639
transform 1 0 0 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 828 0 1 0
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_1
timestamp 1755005639
transform 1 0 828 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_2
timestamp 1755005639
transform 1 0 828 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_3
timestamp 1755005639
transform 1 0 828 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_4
timestamp 1755005639
transform 1 0 828 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_5
timestamp 1755005639
transform 1 0 828 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 736 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1755005639
transform 1 0 736 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 2668 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1755005639
transform 1 0 2668 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1755005639
transform 1 0 2668 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1755005639
transform 1 0 2668 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1755005639
transform 1 0 2668 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1755005639
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
<< labels >>
flabel metal4 20 -48 260 3312 1 FreeSans 160 0 0 0 VDPWR
port 1 n power input
flabel metal4 340 -48 580 3312 1 FreeSans 160 0 0 0 VGND
port 0 n ground input
<< end >>
