magic
tech sky130A
magscale 1 2
timestamp 1756220169
<< nwell >>
rect -2757 -1047 2757 1047
<< mvpmos >>
rect -2499 -750 -2399 750
rect -2341 -750 -2241 750
rect -2183 -750 -2083 750
rect -2025 -750 -1925 750
rect -1867 -750 -1767 750
rect -1709 -750 -1609 750
rect -1551 -750 -1451 750
rect -1393 -750 -1293 750
rect -1235 -750 -1135 750
rect -1077 -750 -977 750
rect -919 -750 -819 750
rect -761 -750 -661 750
rect -603 -750 -503 750
rect -445 -750 -345 750
rect -287 -750 -187 750
rect -129 -750 -29 750
rect 29 -750 129 750
rect 187 -750 287 750
rect 345 -750 445 750
rect 503 -750 603 750
rect 661 -750 761 750
rect 819 -750 919 750
rect 977 -750 1077 750
rect 1135 -750 1235 750
rect 1293 -750 1393 750
rect 1451 -750 1551 750
rect 1609 -750 1709 750
rect 1767 -750 1867 750
rect 1925 -750 2025 750
rect 2083 -750 2183 750
rect 2241 -750 2341 750
rect 2399 -750 2499 750
<< mvpdiff >>
rect -2557 738 -2499 750
rect -2557 -738 -2545 738
rect -2511 -738 -2499 738
rect -2557 -750 -2499 -738
rect -2399 738 -2341 750
rect -2399 -738 -2387 738
rect -2353 -738 -2341 738
rect -2399 -750 -2341 -738
rect -2241 738 -2183 750
rect -2241 -738 -2229 738
rect -2195 -738 -2183 738
rect -2241 -750 -2183 -738
rect -2083 738 -2025 750
rect -2083 -738 -2071 738
rect -2037 -738 -2025 738
rect -2083 -750 -2025 -738
rect -1925 738 -1867 750
rect -1925 -738 -1913 738
rect -1879 -738 -1867 738
rect -1925 -750 -1867 -738
rect -1767 738 -1709 750
rect -1767 -738 -1755 738
rect -1721 -738 -1709 738
rect -1767 -750 -1709 -738
rect -1609 738 -1551 750
rect -1609 -738 -1597 738
rect -1563 -738 -1551 738
rect -1609 -750 -1551 -738
rect -1451 738 -1393 750
rect -1451 -738 -1439 738
rect -1405 -738 -1393 738
rect -1451 -750 -1393 -738
rect -1293 738 -1235 750
rect -1293 -738 -1281 738
rect -1247 -738 -1235 738
rect -1293 -750 -1235 -738
rect -1135 738 -1077 750
rect -1135 -738 -1123 738
rect -1089 -738 -1077 738
rect -1135 -750 -1077 -738
rect -977 738 -919 750
rect -977 -738 -965 738
rect -931 -738 -919 738
rect -977 -750 -919 -738
rect -819 738 -761 750
rect -819 -738 -807 738
rect -773 -738 -761 738
rect -819 -750 -761 -738
rect -661 738 -603 750
rect -661 -738 -649 738
rect -615 -738 -603 738
rect -661 -750 -603 -738
rect -503 738 -445 750
rect -503 -738 -491 738
rect -457 -738 -445 738
rect -503 -750 -445 -738
rect -345 738 -287 750
rect -345 -738 -333 738
rect -299 -738 -287 738
rect -345 -750 -287 -738
rect -187 738 -129 750
rect -187 -738 -175 738
rect -141 -738 -129 738
rect -187 -750 -129 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 129 738 187 750
rect 129 -738 141 738
rect 175 -738 187 738
rect 129 -750 187 -738
rect 287 738 345 750
rect 287 -738 299 738
rect 333 -738 345 738
rect 287 -750 345 -738
rect 445 738 503 750
rect 445 -738 457 738
rect 491 -738 503 738
rect 445 -750 503 -738
rect 603 738 661 750
rect 603 -738 615 738
rect 649 -738 661 738
rect 603 -750 661 -738
rect 761 738 819 750
rect 761 -738 773 738
rect 807 -738 819 738
rect 761 -750 819 -738
rect 919 738 977 750
rect 919 -738 931 738
rect 965 -738 977 738
rect 919 -750 977 -738
rect 1077 738 1135 750
rect 1077 -738 1089 738
rect 1123 -738 1135 738
rect 1077 -750 1135 -738
rect 1235 738 1293 750
rect 1235 -738 1247 738
rect 1281 -738 1293 738
rect 1235 -750 1293 -738
rect 1393 738 1451 750
rect 1393 -738 1405 738
rect 1439 -738 1451 738
rect 1393 -750 1451 -738
rect 1551 738 1609 750
rect 1551 -738 1563 738
rect 1597 -738 1609 738
rect 1551 -750 1609 -738
rect 1709 738 1767 750
rect 1709 -738 1721 738
rect 1755 -738 1767 738
rect 1709 -750 1767 -738
rect 1867 738 1925 750
rect 1867 -738 1879 738
rect 1913 -738 1925 738
rect 1867 -750 1925 -738
rect 2025 738 2083 750
rect 2025 -738 2037 738
rect 2071 -738 2083 738
rect 2025 -750 2083 -738
rect 2183 738 2241 750
rect 2183 -738 2195 738
rect 2229 -738 2241 738
rect 2183 -750 2241 -738
rect 2341 738 2399 750
rect 2341 -738 2353 738
rect 2387 -738 2399 738
rect 2341 -750 2399 -738
rect 2499 738 2557 750
rect 2499 -738 2511 738
rect 2545 -738 2557 738
rect 2499 -750 2557 -738
<< mvpdiffc >>
rect -2545 -738 -2511 738
rect -2387 -738 -2353 738
rect -2229 -738 -2195 738
rect -2071 -738 -2037 738
rect -1913 -738 -1879 738
rect -1755 -738 -1721 738
rect -1597 -738 -1563 738
rect -1439 -738 -1405 738
rect -1281 -738 -1247 738
rect -1123 -738 -1089 738
rect -965 -738 -931 738
rect -807 -738 -773 738
rect -649 -738 -615 738
rect -491 -738 -457 738
rect -333 -738 -299 738
rect -175 -738 -141 738
rect -17 -738 17 738
rect 141 -738 175 738
rect 299 -738 333 738
rect 457 -738 491 738
rect 615 -738 649 738
rect 773 -738 807 738
rect 931 -738 965 738
rect 1089 -738 1123 738
rect 1247 -738 1281 738
rect 1405 -738 1439 738
rect 1563 -738 1597 738
rect 1721 -738 1755 738
rect 1879 -738 1913 738
rect 2037 -738 2071 738
rect 2195 -738 2229 738
rect 2353 -738 2387 738
rect 2511 -738 2545 738
<< mvnsubdiff >>
rect -2691 969 2691 981
rect -2691 935 -2583 969
rect 2583 935 2691 969
rect -2691 923 2691 935
rect -2691 873 -2633 923
rect -2691 -873 -2679 873
rect -2645 -873 -2633 873
rect 2633 873 2691 923
rect -2691 -923 -2633 -873
rect 2633 -873 2645 873
rect 2679 -873 2691 873
rect 2633 -923 2691 -873
rect -2691 -935 2691 -923
rect -2691 -969 -2583 -935
rect 2583 -969 2691 -935
rect -2691 -981 2691 -969
<< mvnsubdiffcont >>
rect -2583 935 2583 969
rect -2679 -873 -2645 873
rect 2645 -873 2679 873
rect -2583 -969 2583 -935
<< poly >>
rect -2499 831 -2399 847
rect -2499 797 -2483 831
rect -2415 797 -2399 831
rect -2499 750 -2399 797
rect -2341 831 -2241 847
rect -2341 797 -2325 831
rect -2257 797 -2241 831
rect -2341 750 -2241 797
rect -2183 831 -2083 847
rect -2183 797 -2167 831
rect -2099 797 -2083 831
rect -2183 750 -2083 797
rect -2025 831 -1925 847
rect -2025 797 -2009 831
rect -1941 797 -1925 831
rect -2025 750 -1925 797
rect -1867 831 -1767 847
rect -1867 797 -1851 831
rect -1783 797 -1767 831
rect -1867 750 -1767 797
rect -1709 831 -1609 847
rect -1709 797 -1693 831
rect -1625 797 -1609 831
rect -1709 750 -1609 797
rect -1551 831 -1451 847
rect -1551 797 -1535 831
rect -1467 797 -1451 831
rect -1551 750 -1451 797
rect -1393 831 -1293 847
rect -1393 797 -1377 831
rect -1309 797 -1293 831
rect -1393 750 -1293 797
rect -1235 831 -1135 847
rect -1235 797 -1219 831
rect -1151 797 -1135 831
rect -1235 750 -1135 797
rect -1077 831 -977 847
rect -1077 797 -1061 831
rect -993 797 -977 831
rect -1077 750 -977 797
rect -919 831 -819 847
rect -919 797 -903 831
rect -835 797 -819 831
rect -919 750 -819 797
rect -761 831 -661 847
rect -761 797 -745 831
rect -677 797 -661 831
rect -761 750 -661 797
rect -603 831 -503 847
rect -603 797 -587 831
rect -519 797 -503 831
rect -603 750 -503 797
rect -445 831 -345 847
rect -445 797 -429 831
rect -361 797 -345 831
rect -445 750 -345 797
rect -287 831 -187 847
rect -287 797 -271 831
rect -203 797 -187 831
rect -287 750 -187 797
rect -129 831 -29 847
rect -129 797 -113 831
rect -45 797 -29 831
rect -129 750 -29 797
rect 29 831 129 847
rect 29 797 45 831
rect 113 797 129 831
rect 29 750 129 797
rect 187 831 287 847
rect 187 797 203 831
rect 271 797 287 831
rect 187 750 287 797
rect 345 831 445 847
rect 345 797 361 831
rect 429 797 445 831
rect 345 750 445 797
rect 503 831 603 847
rect 503 797 519 831
rect 587 797 603 831
rect 503 750 603 797
rect 661 831 761 847
rect 661 797 677 831
rect 745 797 761 831
rect 661 750 761 797
rect 819 831 919 847
rect 819 797 835 831
rect 903 797 919 831
rect 819 750 919 797
rect 977 831 1077 847
rect 977 797 993 831
rect 1061 797 1077 831
rect 977 750 1077 797
rect 1135 831 1235 847
rect 1135 797 1151 831
rect 1219 797 1235 831
rect 1135 750 1235 797
rect 1293 831 1393 847
rect 1293 797 1309 831
rect 1377 797 1393 831
rect 1293 750 1393 797
rect 1451 831 1551 847
rect 1451 797 1467 831
rect 1535 797 1551 831
rect 1451 750 1551 797
rect 1609 831 1709 847
rect 1609 797 1625 831
rect 1693 797 1709 831
rect 1609 750 1709 797
rect 1767 831 1867 847
rect 1767 797 1783 831
rect 1851 797 1867 831
rect 1767 750 1867 797
rect 1925 831 2025 847
rect 1925 797 1941 831
rect 2009 797 2025 831
rect 1925 750 2025 797
rect 2083 831 2183 847
rect 2083 797 2099 831
rect 2167 797 2183 831
rect 2083 750 2183 797
rect 2241 831 2341 847
rect 2241 797 2257 831
rect 2325 797 2341 831
rect 2241 750 2341 797
rect 2399 831 2499 847
rect 2399 797 2415 831
rect 2483 797 2499 831
rect 2399 750 2499 797
rect -2499 -797 -2399 -750
rect -2499 -831 -2483 -797
rect -2415 -831 -2399 -797
rect -2499 -847 -2399 -831
rect -2341 -797 -2241 -750
rect -2341 -831 -2325 -797
rect -2257 -831 -2241 -797
rect -2341 -847 -2241 -831
rect -2183 -797 -2083 -750
rect -2183 -831 -2167 -797
rect -2099 -831 -2083 -797
rect -2183 -847 -2083 -831
rect -2025 -797 -1925 -750
rect -2025 -831 -2009 -797
rect -1941 -831 -1925 -797
rect -2025 -847 -1925 -831
rect -1867 -797 -1767 -750
rect -1867 -831 -1851 -797
rect -1783 -831 -1767 -797
rect -1867 -847 -1767 -831
rect -1709 -797 -1609 -750
rect -1709 -831 -1693 -797
rect -1625 -831 -1609 -797
rect -1709 -847 -1609 -831
rect -1551 -797 -1451 -750
rect -1551 -831 -1535 -797
rect -1467 -831 -1451 -797
rect -1551 -847 -1451 -831
rect -1393 -797 -1293 -750
rect -1393 -831 -1377 -797
rect -1309 -831 -1293 -797
rect -1393 -847 -1293 -831
rect -1235 -797 -1135 -750
rect -1235 -831 -1219 -797
rect -1151 -831 -1135 -797
rect -1235 -847 -1135 -831
rect -1077 -797 -977 -750
rect -1077 -831 -1061 -797
rect -993 -831 -977 -797
rect -1077 -847 -977 -831
rect -919 -797 -819 -750
rect -919 -831 -903 -797
rect -835 -831 -819 -797
rect -919 -847 -819 -831
rect -761 -797 -661 -750
rect -761 -831 -745 -797
rect -677 -831 -661 -797
rect -761 -847 -661 -831
rect -603 -797 -503 -750
rect -603 -831 -587 -797
rect -519 -831 -503 -797
rect -603 -847 -503 -831
rect -445 -797 -345 -750
rect -445 -831 -429 -797
rect -361 -831 -345 -797
rect -445 -847 -345 -831
rect -287 -797 -187 -750
rect -287 -831 -271 -797
rect -203 -831 -187 -797
rect -287 -847 -187 -831
rect -129 -797 -29 -750
rect -129 -831 -113 -797
rect -45 -831 -29 -797
rect -129 -847 -29 -831
rect 29 -797 129 -750
rect 29 -831 45 -797
rect 113 -831 129 -797
rect 29 -847 129 -831
rect 187 -797 287 -750
rect 187 -831 203 -797
rect 271 -831 287 -797
rect 187 -847 287 -831
rect 345 -797 445 -750
rect 345 -831 361 -797
rect 429 -831 445 -797
rect 345 -847 445 -831
rect 503 -797 603 -750
rect 503 -831 519 -797
rect 587 -831 603 -797
rect 503 -847 603 -831
rect 661 -797 761 -750
rect 661 -831 677 -797
rect 745 -831 761 -797
rect 661 -847 761 -831
rect 819 -797 919 -750
rect 819 -831 835 -797
rect 903 -831 919 -797
rect 819 -847 919 -831
rect 977 -797 1077 -750
rect 977 -831 993 -797
rect 1061 -831 1077 -797
rect 977 -847 1077 -831
rect 1135 -797 1235 -750
rect 1135 -831 1151 -797
rect 1219 -831 1235 -797
rect 1135 -847 1235 -831
rect 1293 -797 1393 -750
rect 1293 -831 1309 -797
rect 1377 -831 1393 -797
rect 1293 -847 1393 -831
rect 1451 -797 1551 -750
rect 1451 -831 1467 -797
rect 1535 -831 1551 -797
rect 1451 -847 1551 -831
rect 1609 -797 1709 -750
rect 1609 -831 1625 -797
rect 1693 -831 1709 -797
rect 1609 -847 1709 -831
rect 1767 -797 1867 -750
rect 1767 -831 1783 -797
rect 1851 -831 1867 -797
rect 1767 -847 1867 -831
rect 1925 -797 2025 -750
rect 1925 -831 1941 -797
rect 2009 -831 2025 -797
rect 1925 -847 2025 -831
rect 2083 -797 2183 -750
rect 2083 -831 2099 -797
rect 2167 -831 2183 -797
rect 2083 -847 2183 -831
rect 2241 -797 2341 -750
rect 2241 -831 2257 -797
rect 2325 -831 2341 -797
rect 2241 -847 2341 -831
rect 2399 -797 2499 -750
rect 2399 -831 2415 -797
rect 2483 -831 2499 -797
rect 2399 -847 2499 -831
<< polycont >>
rect -2483 797 -2415 831
rect -2325 797 -2257 831
rect -2167 797 -2099 831
rect -2009 797 -1941 831
rect -1851 797 -1783 831
rect -1693 797 -1625 831
rect -1535 797 -1467 831
rect -1377 797 -1309 831
rect -1219 797 -1151 831
rect -1061 797 -993 831
rect -903 797 -835 831
rect -745 797 -677 831
rect -587 797 -519 831
rect -429 797 -361 831
rect -271 797 -203 831
rect -113 797 -45 831
rect 45 797 113 831
rect 203 797 271 831
rect 361 797 429 831
rect 519 797 587 831
rect 677 797 745 831
rect 835 797 903 831
rect 993 797 1061 831
rect 1151 797 1219 831
rect 1309 797 1377 831
rect 1467 797 1535 831
rect 1625 797 1693 831
rect 1783 797 1851 831
rect 1941 797 2009 831
rect 2099 797 2167 831
rect 2257 797 2325 831
rect 2415 797 2483 831
rect -2483 -831 -2415 -797
rect -2325 -831 -2257 -797
rect -2167 -831 -2099 -797
rect -2009 -831 -1941 -797
rect -1851 -831 -1783 -797
rect -1693 -831 -1625 -797
rect -1535 -831 -1467 -797
rect -1377 -831 -1309 -797
rect -1219 -831 -1151 -797
rect -1061 -831 -993 -797
rect -903 -831 -835 -797
rect -745 -831 -677 -797
rect -587 -831 -519 -797
rect -429 -831 -361 -797
rect -271 -831 -203 -797
rect -113 -831 -45 -797
rect 45 -831 113 -797
rect 203 -831 271 -797
rect 361 -831 429 -797
rect 519 -831 587 -797
rect 677 -831 745 -797
rect 835 -831 903 -797
rect 993 -831 1061 -797
rect 1151 -831 1219 -797
rect 1309 -831 1377 -797
rect 1467 -831 1535 -797
rect 1625 -831 1693 -797
rect 1783 -831 1851 -797
rect 1941 -831 2009 -797
rect 2099 -831 2167 -797
rect 2257 -831 2325 -797
rect 2415 -831 2483 -797
<< locali >>
rect -2679 935 -2583 969
rect 2583 935 2679 969
rect -2679 873 -2645 935
rect 2645 873 2679 935
rect -2499 797 -2483 831
rect -2415 797 -2399 831
rect -2341 797 -2325 831
rect -2257 797 -2241 831
rect -2183 797 -2167 831
rect -2099 797 -2083 831
rect -2025 797 -2009 831
rect -1941 797 -1925 831
rect -1867 797 -1851 831
rect -1783 797 -1767 831
rect -1709 797 -1693 831
rect -1625 797 -1609 831
rect -1551 797 -1535 831
rect -1467 797 -1451 831
rect -1393 797 -1377 831
rect -1309 797 -1293 831
rect -1235 797 -1219 831
rect -1151 797 -1135 831
rect -1077 797 -1061 831
rect -993 797 -977 831
rect -919 797 -903 831
rect -835 797 -819 831
rect -761 797 -745 831
rect -677 797 -661 831
rect -603 797 -587 831
rect -519 797 -503 831
rect -445 797 -429 831
rect -361 797 -345 831
rect -287 797 -271 831
rect -203 797 -187 831
rect -129 797 -113 831
rect -45 797 -29 831
rect 29 797 45 831
rect 113 797 129 831
rect 187 797 203 831
rect 271 797 287 831
rect 345 797 361 831
rect 429 797 445 831
rect 503 797 519 831
rect 587 797 603 831
rect 661 797 677 831
rect 745 797 761 831
rect 819 797 835 831
rect 903 797 919 831
rect 977 797 993 831
rect 1061 797 1077 831
rect 1135 797 1151 831
rect 1219 797 1235 831
rect 1293 797 1309 831
rect 1377 797 1393 831
rect 1451 797 1467 831
rect 1535 797 1551 831
rect 1609 797 1625 831
rect 1693 797 1709 831
rect 1767 797 1783 831
rect 1851 797 1867 831
rect 1925 797 1941 831
rect 2009 797 2025 831
rect 2083 797 2099 831
rect 2167 797 2183 831
rect 2241 797 2257 831
rect 2325 797 2341 831
rect 2399 797 2415 831
rect 2483 797 2499 831
rect -2545 738 -2511 754
rect -2545 -754 -2511 -738
rect -2387 738 -2353 754
rect -2387 -754 -2353 -738
rect -2229 738 -2195 754
rect -2229 -754 -2195 -738
rect -2071 738 -2037 754
rect -2071 -754 -2037 -738
rect -1913 738 -1879 754
rect -1913 -754 -1879 -738
rect -1755 738 -1721 754
rect -1755 -754 -1721 -738
rect -1597 738 -1563 754
rect -1597 -754 -1563 -738
rect -1439 738 -1405 754
rect -1439 -754 -1405 -738
rect -1281 738 -1247 754
rect -1281 -754 -1247 -738
rect -1123 738 -1089 754
rect -1123 -754 -1089 -738
rect -965 738 -931 754
rect -965 -754 -931 -738
rect -807 738 -773 754
rect -807 -754 -773 -738
rect -649 738 -615 754
rect -649 -754 -615 -738
rect -491 738 -457 754
rect -491 -754 -457 -738
rect -333 738 -299 754
rect -333 -754 -299 -738
rect -175 738 -141 754
rect -175 -754 -141 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 141 738 175 754
rect 141 -754 175 -738
rect 299 738 333 754
rect 299 -754 333 -738
rect 457 738 491 754
rect 457 -754 491 -738
rect 615 738 649 754
rect 615 -754 649 -738
rect 773 738 807 754
rect 773 -754 807 -738
rect 931 738 965 754
rect 931 -754 965 -738
rect 1089 738 1123 754
rect 1089 -754 1123 -738
rect 1247 738 1281 754
rect 1247 -754 1281 -738
rect 1405 738 1439 754
rect 1405 -754 1439 -738
rect 1563 738 1597 754
rect 1563 -754 1597 -738
rect 1721 738 1755 754
rect 1721 -754 1755 -738
rect 1879 738 1913 754
rect 1879 -754 1913 -738
rect 2037 738 2071 754
rect 2037 -754 2071 -738
rect 2195 738 2229 754
rect 2195 -754 2229 -738
rect 2353 738 2387 754
rect 2353 -754 2387 -738
rect 2511 738 2545 754
rect 2511 -754 2545 -738
rect -2499 -831 -2483 -797
rect -2415 -831 -2399 -797
rect -2341 -831 -2325 -797
rect -2257 -831 -2241 -797
rect -2183 -831 -2167 -797
rect -2099 -831 -2083 -797
rect -2025 -831 -2009 -797
rect -1941 -831 -1925 -797
rect -1867 -831 -1851 -797
rect -1783 -831 -1767 -797
rect -1709 -831 -1693 -797
rect -1625 -831 -1609 -797
rect -1551 -831 -1535 -797
rect -1467 -831 -1451 -797
rect -1393 -831 -1377 -797
rect -1309 -831 -1293 -797
rect -1235 -831 -1219 -797
rect -1151 -831 -1135 -797
rect -1077 -831 -1061 -797
rect -993 -831 -977 -797
rect -919 -831 -903 -797
rect -835 -831 -819 -797
rect -761 -831 -745 -797
rect -677 -831 -661 -797
rect -603 -831 -587 -797
rect -519 -831 -503 -797
rect -445 -831 -429 -797
rect -361 -831 -345 -797
rect -287 -831 -271 -797
rect -203 -831 -187 -797
rect -129 -831 -113 -797
rect -45 -831 -29 -797
rect 29 -831 45 -797
rect 113 -831 129 -797
rect 187 -831 203 -797
rect 271 -831 287 -797
rect 345 -831 361 -797
rect 429 -831 445 -797
rect 503 -831 519 -797
rect 587 -831 603 -797
rect 661 -831 677 -797
rect 745 -831 761 -797
rect 819 -831 835 -797
rect 903 -831 919 -797
rect 977 -831 993 -797
rect 1061 -831 1077 -797
rect 1135 -831 1151 -797
rect 1219 -831 1235 -797
rect 1293 -831 1309 -797
rect 1377 -831 1393 -797
rect 1451 -831 1467 -797
rect 1535 -831 1551 -797
rect 1609 -831 1625 -797
rect 1693 -831 1709 -797
rect 1767 -831 1783 -797
rect 1851 -831 1867 -797
rect 1925 -831 1941 -797
rect 2009 -831 2025 -797
rect 2083 -831 2099 -797
rect 2167 -831 2183 -797
rect 2241 -831 2257 -797
rect 2325 -831 2341 -797
rect 2399 -831 2415 -797
rect 2483 -831 2499 -797
rect -2679 -935 -2645 -873
rect 2645 -935 2679 -873
rect -2679 -969 -2583 -935
rect 2583 -969 2679 -935
<< viali >>
rect -2483 797 -2415 831
rect -2325 797 -2257 831
rect -2167 797 -2099 831
rect -2009 797 -1941 831
rect -1851 797 -1783 831
rect -1693 797 -1625 831
rect -1535 797 -1467 831
rect -1377 797 -1309 831
rect -1219 797 -1151 831
rect -1061 797 -993 831
rect -903 797 -835 831
rect -745 797 -677 831
rect -587 797 -519 831
rect -429 797 -361 831
rect -271 797 -203 831
rect -113 797 -45 831
rect 45 797 113 831
rect 203 797 271 831
rect 361 797 429 831
rect 519 797 587 831
rect 677 797 745 831
rect 835 797 903 831
rect 993 797 1061 831
rect 1151 797 1219 831
rect 1309 797 1377 831
rect 1467 797 1535 831
rect 1625 797 1693 831
rect 1783 797 1851 831
rect 1941 797 2009 831
rect 2099 797 2167 831
rect 2257 797 2325 831
rect 2415 797 2483 831
rect -2545 -738 -2511 738
rect -2387 -738 -2353 738
rect -2229 -738 -2195 738
rect -2071 -738 -2037 738
rect -1913 -738 -1879 738
rect -1755 -738 -1721 738
rect -1597 -738 -1563 738
rect -1439 -738 -1405 738
rect -1281 -738 -1247 738
rect -1123 -738 -1089 738
rect -965 -738 -931 738
rect -807 -738 -773 738
rect -649 -738 -615 738
rect -491 -738 -457 738
rect -333 -738 -299 738
rect -175 -738 -141 738
rect -17 -738 17 738
rect 141 -738 175 738
rect 299 -738 333 738
rect 457 -738 491 738
rect 615 -738 649 738
rect 773 -738 807 738
rect 931 -738 965 738
rect 1089 -738 1123 738
rect 1247 -738 1281 738
rect 1405 -738 1439 738
rect 1563 -738 1597 738
rect 1721 -738 1755 738
rect 1879 -738 1913 738
rect 2037 -738 2071 738
rect 2195 -738 2229 738
rect 2353 -738 2387 738
rect 2511 -738 2545 738
rect -2483 -831 -2415 -797
rect -2325 -831 -2257 -797
rect -2167 -831 -2099 -797
rect -2009 -831 -1941 -797
rect -1851 -831 -1783 -797
rect -1693 -831 -1625 -797
rect -1535 -831 -1467 -797
rect -1377 -831 -1309 -797
rect -1219 -831 -1151 -797
rect -1061 -831 -993 -797
rect -903 -831 -835 -797
rect -745 -831 -677 -797
rect -587 -831 -519 -797
rect -429 -831 -361 -797
rect -271 -831 -203 -797
rect -113 -831 -45 -797
rect 45 -831 113 -797
rect 203 -831 271 -797
rect 361 -831 429 -797
rect 519 -831 587 -797
rect 677 -831 745 -797
rect 835 -831 903 -797
rect 993 -831 1061 -797
rect 1151 -831 1219 -797
rect 1309 -831 1377 -797
rect 1467 -831 1535 -797
rect 1625 -831 1693 -797
rect 1783 -831 1851 -797
rect 1941 -831 2009 -797
rect 2099 -831 2167 -797
rect 2257 -831 2325 -797
rect 2415 -831 2483 -797
<< metal1 >>
rect -2495 831 -2403 837
rect -2495 797 -2483 831
rect -2415 797 -2403 831
rect -2495 791 -2403 797
rect -2337 831 -2245 837
rect -2337 797 -2325 831
rect -2257 797 -2245 831
rect -2337 791 -2245 797
rect -2179 831 -2087 837
rect -2179 797 -2167 831
rect -2099 797 -2087 831
rect -2179 791 -2087 797
rect -2021 831 -1929 837
rect -2021 797 -2009 831
rect -1941 797 -1929 831
rect -2021 791 -1929 797
rect -1863 831 -1771 837
rect -1863 797 -1851 831
rect -1783 797 -1771 831
rect -1863 791 -1771 797
rect -1705 831 -1613 837
rect -1705 797 -1693 831
rect -1625 797 -1613 831
rect -1705 791 -1613 797
rect -1547 831 -1455 837
rect -1547 797 -1535 831
rect -1467 797 -1455 831
rect -1547 791 -1455 797
rect -1389 831 -1297 837
rect -1389 797 -1377 831
rect -1309 797 -1297 831
rect -1389 791 -1297 797
rect -1231 831 -1139 837
rect -1231 797 -1219 831
rect -1151 797 -1139 831
rect -1231 791 -1139 797
rect -1073 831 -981 837
rect -1073 797 -1061 831
rect -993 797 -981 831
rect -1073 791 -981 797
rect -915 831 -823 837
rect -915 797 -903 831
rect -835 797 -823 831
rect -915 791 -823 797
rect -757 831 -665 837
rect -757 797 -745 831
rect -677 797 -665 831
rect -757 791 -665 797
rect -599 831 -507 837
rect -599 797 -587 831
rect -519 797 -507 831
rect -599 791 -507 797
rect -441 831 -349 837
rect -441 797 -429 831
rect -361 797 -349 831
rect -441 791 -349 797
rect -283 831 -191 837
rect -283 797 -271 831
rect -203 797 -191 831
rect -283 791 -191 797
rect -125 831 -33 837
rect -125 797 -113 831
rect -45 797 -33 831
rect -125 791 -33 797
rect 33 831 125 837
rect 33 797 45 831
rect 113 797 125 831
rect 33 791 125 797
rect 191 831 283 837
rect 191 797 203 831
rect 271 797 283 831
rect 191 791 283 797
rect 349 831 441 837
rect 349 797 361 831
rect 429 797 441 831
rect 349 791 441 797
rect 507 831 599 837
rect 507 797 519 831
rect 587 797 599 831
rect 507 791 599 797
rect 665 831 757 837
rect 665 797 677 831
rect 745 797 757 831
rect 665 791 757 797
rect 823 831 915 837
rect 823 797 835 831
rect 903 797 915 831
rect 823 791 915 797
rect 981 831 1073 837
rect 981 797 993 831
rect 1061 797 1073 831
rect 981 791 1073 797
rect 1139 831 1231 837
rect 1139 797 1151 831
rect 1219 797 1231 831
rect 1139 791 1231 797
rect 1297 831 1389 837
rect 1297 797 1309 831
rect 1377 797 1389 831
rect 1297 791 1389 797
rect 1455 831 1547 837
rect 1455 797 1467 831
rect 1535 797 1547 831
rect 1455 791 1547 797
rect 1613 831 1705 837
rect 1613 797 1625 831
rect 1693 797 1705 831
rect 1613 791 1705 797
rect 1771 831 1863 837
rect 1771 797 1783 831
rect 1851 797 1863 831
rect 1771 791 1863 797
rect 1929 831 2021 837
rect 1929 797 1941 831
rect 2009 797 2021 831
rect 1929 791 2021 797
rect 2087 831 2179 837
rect 2087 797 2099 831
rect 2167 797 2179 831
rect 2087 791 2179 797
rect 2245 831 2337 837
rect 2245 797 2257 831
rect 2325 797 2337 831
rect 2245 791 2337 797
rect 2403 831 2495 837
rect 2403 797 2415 831
rect 2483 797 2495 831
rect 2403 791 2495 797
rect -2551 738 -2505 750
rect -2551 -738 -2545 738
rect -2511 -738 -2505 738
rect -2551 -750 -2505 -738
rect -2393 738 -2347 750
rect -2393 -738 -2387 738
rect -2353 -738 -2347 738
rect -2393 -750 -2347 -738
rect -2235 738 -2189 750
rect -2235 -738 -2229 738
rect -2195 -738 -2189 738
rect -2235 -750 -2189 -738
rect -2077 738 -2031 750
rect -2077 -738 -2071 738
rect -2037 -738 -2031 738
rect -2077 -750 -2031 -738
rect -1919 738 -1873 750
rect -1919 -738 -1913 738
rect -1879 -738 -1873 738
rect -1919 -750 -1873 -738
rect -1761 738 -1715 750
rect -1761 -738 -1755 738
rect -1721 -738 -1715 738
rect -1761 -750 -1715 -738
rect -1603 738 -1557 750
rect -1603 -738 -1597 738
rect -1563 -738 -1557 738
rect -1603 -750 -1557 -738
rect -1445 738 -1399 750
rect -1445 -738 -1439 738
rect -1405 -738 -1399 738
rect -1445 -750 -1399 -738
rect -1287 738 -1241 750
rect -1287 -738 -1281 738
rect -1247 -738 -1241 738
rect -1287 -750 -1241 -738
rect -1129 738 -1083 750
rect -1129 -738 -1123 738
rect -1089 -738 -1083 738
rect -1129 -750 -1083 -738
rect -971 738 -925 750
rect -971 -738 -965 738
rect -931 -738 -925 738
rect -971 -750 -925 -738
rect -813 738 -767 750
rect -813 -738 -807 738
rect -773 -738 -767 738
rect -813 -750 -767 -738
rect -655 738 -609 750
rect -655 -738 -649 738
rect -615 -738 -609 738
rect -655 -750 -609 -738
rect -497 738 -451 750
rect -497 -738 -491 738
rect -457 -738 -451 738
rect -497 -750 -451 -738
rect -339 738 -293 750
rect -339 -738 -333 738
rect -299 -738 -293 738
rect -339 -750 -293 -738
rect -181 738 -135 750
rect -181 -738 -175 738
rect -141 -738 -135 738
rect -181 -750 -135 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 135 738 181 750
rect 135 -738 141 738
rect 175 -738 181 738
rect 135 -750 181 -738
rect 293 738 339 750
rect 293 -738 299 738
rect 333 -738 339 738
rect 293 -750 339 -738
rect 451 738 497 750
rect 451 -738 457 738
rect 491 -738 497 738
rect 451 -750 497 -738
rect 609 738 655 750
rect 609 -738 615 738
rect 649 -738 655 738
rect 609 -750 655 -738
rect 767 738 813 750
rect 767 -738 773 738
rect 807 -738 813 738
rect 767 -750 813 -738
rect 925 738 971 750
rect 925 -738 931 738
rect 965 -738 971 738
rect 925 -750 971 -738
rect 1083 738 1129 750
rect 1083 -738 1089 738
rect 1123 -738 1129 738
rect 1083 -750 1129 -738
rect 1241 738 1287 750
rect 1241 -738 1247 738
rect 1281 -738 1287 738
rect 1241 -750 1287 -738
rect 1399 738 1445 750
rect 1399 -738 1405 738
rect 1439 -738 1445 738
rect 1399 -750 1445 -738
rect 1557 738 1603 750
rect 1557 -738 1563 738
rect 1597 -738 1603 738
rect 1557 -750 1603 -738
rect 1715 738 1761 750
rect 1715 -738 1721 738
rect 1755 -738 1761 738
rect 1715 -750 1761 -738
rect 1873 738 1919 750
rect 1873 -738 1879 738
rect 1913 -738 1919 738
rect 1873 -750 1919 -738
rect 2031 738 2077 750
rect 2031 -738 2037 738
rect 2071 -738 2077 738
rect 2031 -750 2077 -738
rect 2189 738 2235 750
rect 2189 -738 2195 738
rect 2229 -738 2235 738
rect 2189 -750 2235 -738
rect 2347 738 2393 750
rect 2347 -738 2353 738
rect 2387 -738 2393 738
rect 2347 -750 2393 -738
rect 2505 738 2551 750
rect 2505 -738 2511 738
rect 2545 -738 2551 738
rect 2505 -750 2551 -738
rect -2495 -797 -2403 -791
rect -2495 -831 -2483 -797
rect -2415 -831 -2403 -797
rect -2495 -837 -2403 -831
rect -2337 -797 -2245 -791
rect -2337 -831 -2325 -797
rect -2257 -831 -2245 -797
rect -2337 -837 -2245 -831
rect -2179 -797 -2087 -791
rect -2179 -831 -2167 -797
rect -2099 -831 -2087 -797
rect -2179 -837 -2087 -831
rect -2021 -797 -1929 -791
rect -2021 -831 -2009 -797
rect -1941 -831 -1929 -797
rect -2021 -837 -1929 -831
rect -1863 -797 -1771 -791
rect -1863 -831 -1851 -797
rect -1783 -831 -1771 -797
rect -1863 -837 -1771 -831
rect -1705 -797 -1613 -791
rect -1705 -831 -1693 -797
rect -1625 -831 -1613 -797
rect -1705 -837 -1613 -831
rect -1547 -797 -1455 -791
rect -1547 -831 -1535 -797
rect -1467 -831 -1455 -797
rect -1547 -837 -1455 -831
rect -1389 -797 -1297 -791
rect -1389 -831 -1377 -797
rect -1309 -831 -1297 -797
rect -1389 -837 -1297 -831
rect -1231 -797 -1139 -791
rect -1231 -831 -1219 -797
rect -1151 -831 -1139 -797
rect -1231 -837 -1139 -831
rect -1073 -797 -981 -791
rect -1073 -831 -1061 -797
rect -993 -831 -981 -797
rect -1073 -837 -981 -831
rect -915 -797 -823 -791
rect -915 -831 -903 -797
rect -835 -831 -823 -797
rect -915 -837 -823 -831
rect -757 -797 -665 -791
rect -757 -831 -745 -797
rect -677 -831 -665 -797
rect -757 -837 -665 -831
rect -599 -797 -507 -791
rect -599 -831 -587 -797
rect -519 -831 -507 -797
rect -599 -837 -507 -831
rect -441 -797 -349 -791
rect -441 -831 -429 -797
rect -361 -831 -349 -797
rect -441 -837 -349 -831
rect -283 -797 -191 -791
rect -283 -831 -271 -797
rect -203 -831 -191 -797
rect -283 -837 -191 -831
rect -125 -797 -33 -791
rect -125 -831 -113 -797
rect -45 -831 -33 -797
rect -125 -837 -33 -831
rect 33 -797 125 -791
rect 33 -831 45 -797
rect 113 -831 125 -797
rect 33 -837 125 -831
rect 191 -797 283 -791
rect 191 -831 203 -797
rect 271 -831 283 -797
rect 191 -837 283 -831
rect 349 -797 441 -791
rect 349 -831 361 -797
rect 429 -831 441 -797
rect 349 -837 441 -831
rect 507 -797 599 -791
rect 507 -831 519 -797
rect 587 -831 599 -797
rect 507 -837 599 -831
rect 665 -797 757 -791
rect 665 -831 677 -797
rect 745 -831 757 -797
rect 665 -837 757 -831
rect 823 -797 915 -791
rect 823 -831 835 -797
rect 903 -831 915 -797
rect 823 -837 915 -831
rect 981 -797 1073 -791
rect 981 -831 993 -797
rect 1061 -831 1073 -797
rect 981 -837 1073 -831
rect 1139 -797 1231 -791
rect 1139 -831 1151 -797
rect 1219 -831 1231 -797
rect 1139 -837 1231 -831
rect 1297 -797 1389 -791
rect 1297 -831 1309 -797
rect 1377 -831 1389 -797
rect 1297 -837 1389 -831
rect 1455 -797 1547 -791
rect 1455 -831 1467 -797
rect 1535 -831 1547 -797
rect 1455 -837 1547 -831
rect 1613 -797 1705 -791
rect 1613 -831 1625 -797
rect 1693 -831 1705 -797
rect 1613 -837 1705 -831
rect 1771 -797 1863 -791
rect 1771 -831 1783 -797
rect 1851 -831 1863 -797
rect 1771 -837 1863 -831
rect 1929 -797 2021 -791
rect 1929 -831 1941 -797
rect 2009 -831 2021 -797
rect 1929 -837 2021 -831
rect 2087 -797 2179 -791
rect 2087 -831 2099 -797
rect 2167 -831 2179 -797
rect 2087 -837 2179 -831
rect 2245 -797 2337 -791
rect 2245 -831 2257 -797
rect 2325 -831 2337 -797
rect 2245 -837 2337 -831
rect 2403 -797 2495 -791
rect 2403 -831 2415 -797
rect 2483 -831 2495 -797
rect 2403 -837 2495 -831
<< labels >>
rlabel mvnsubdiffcont 0 -952 0 -952 0 B
port 1 nsew
rlabel mvpdiffc -2528 0 -2528 0 0 D0
port 2 nsew
rlabel polycont -2449 814 -2449 814 0 G0
port 3 nsew
rlabel mvpdiffc -2370 0 -2370 0 0 S1
port 4 nsew
rlabel polycont -2291 814 -2291 814 0 G1
port 5 nsew
rlabel mvpdiffc -2212 0 -2212 0 0 D2
port 6 nsew
rlabel polycont -2133 814 -2133 814 0 G2
port 7 nsew
rlabel mvpdiffc -2054 0 -2054 0 0 S3
port 8 nsew
rlabel polycont -1975 814 -1975 814 0 G3
port 9 nsew
rlabel mvpdiffc -1896 0 -1896 0 0 D4
port 10 nsew
rlabel polycont -1817 814 -1817 814 0 G4
port 11 nsew
rlabel mvpdiffc -1738 0 -1738 0 0 S5
port 12 nsew
rlabel polycont -1659 814 -1659 814 0 G5
port 13 nsew
rlabel mvpdiffc -1580 0 -1580 0 0 D6
port 14 nsew
rlabel polycont -1501 814 -1501 814 0 G6
port 15 nsew
rlabel mvpdiffc -1422 0 -1422 0 0 S7
port 16 nsew
rlabel polycont -1343 814 -1343 814 0 G7
port 17 nsew
rlabel mvpdiffc -1264 0 -1264 0 0 D8
port 18 nsew
rlabel polycont -1185 814 -1185 814 0 G8
port 19 nsew
rlabel mvpdiffc -1106 0 -1106 0 0 S9
port 20 nsew
rlabel polycont -1027 814 -1027 814 0 G9
port 21 nsew
rlabel mvpdiffc -948 0 -948 0 0 D10
port 22 nsew
rlabel polycont -869 814 -869 814 0 G10
port 23 nsew
rlabel mvpdiffc -790 0 -790 0 0 S11
port 24 nsew
rlabel polycont -711 814 -711 814 0 G11
port 25 nsew
rlabel mvpdiffc -632 0 -632 0 0 D12
port 26 nsew
rlabel polycont -553 814 -553 814 0 G12
port 27 nsew
rlabel mvpdiffc -474 0 -474 0 0 S13
port 28 nsew
rlabel polycont -395 814 -395 814 0 G13
port 29 nsew
rlabel mvpdiffc -316 0 -316 0 0 D14
port 30 nsew
rlabel polycont -237 814 -237 814 0 G14
port 31 nsew
rlabel mvpdiffc -158 0 -158 0 0 S15
port 32 nsew
rlabel polycont -79 814 -79 814 0 G15
port 33 nsew
rlabel mvpdiffc 0 0 0 0 0 D16
port 34 nsew
rlabel polycont 79 814 79 814 0 G16
port 35 nsew
rlabel mvpdiffc 158 0 158 0 0 S17
port 36 nsew
rlabel polycont 237 814 237 814 0 G17
port 37 nsew
rlabel mvpdiffc 316 0 316 0 0 D18
port 38 nsew
rlabel polycont 395 814 395 814 0 G18
port 39 nsew
rlabel mvpdiffc 474 0 474 0 0 S19
port 40 nsew
rlabel polycont 553 814 553 814 0 G19
port 41 nsew
rlabel mvpdiffc 632 0 632 0 0 D20
port 42 nsew
rlabel polycont 711 814 711 814 0 G20
port 43 nsew
rlabel mvpdiffc 790 0 790 0 0 S21
port 44 nsew
rlabel polycont 869 814 869 814 0 G21
port 45 nsew
rlabel mvpdiffc 948 0 948 0 0 D22
port 46 nsew
rlabel polycont 1027 814 1027 814 0 G22
port 47 nsew
rlabel mvpdiffc 1106 0 1106 0 0 S23
port 48 nsew
rlabel polycont 1185 814 1185 814 0 G23
port 49 nsew
rlabel mvpdiffc 1264 0 1264 0 0 D24
port 50 nsew
rlabel polycont 1343 814 1343 814 0 G24
port 51 nsew
rlabel mvpdiffc 1422 0 1422 0 0 S25
port 52 nsew
rlabel polycont 1501 814 1501 814 0 G25
port 53 nsew
rlabel mvpdiffc 1580 0 1580 0 0 D26
port 54 nsew
rlabel polycont 1659 814 1659 814 0 G26
port 55 nsew
rlabel mvpdiffc 1738 0 1738 0 0 S27
port 56 nsew
rlabel polycont 1817 814 1817 814 0 G27
port 57 nsew
rlabel mvpdiffc 1896 0 1896 0 0 D28
port 58 nsew
rlabel polycont 1975 814 1975 814 0 G28
port 59 nsew
rlabel mvpdiffc 2054 0 2054 0 0 S29
port 60 nsew
rlabel polycont 2133 814 2133 814 0 G29
port 61 nsew
rlabel mvpdiffc 2212 0 2212 0 0 D30
port 62 nsew
rlabel polycont 2291 814 2291 814 0 G30
port 63 nsew
rlabel mvpdiffc 2370 0 2370 0 0 S31
port 64 nsew
rlabel polycont 2449 814 2449 814 0 G31
port 65 nsew
<< properties >>
string FIXED_BBOX -2662 -952 2662 952
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 0.50 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
