magic
tech sky130A
magscale 1 2
timestamp 1756676326
<< viali >>
rect 377 12534 18023 12568
rect 277 10730 311 12468
rect 18089 10730 18123 12468
rect 377 10630 18023 10664
<< metal1 >>
rect 654 12574 660 12577
rect 271 12568 660 12574
rect 712 12574 718 12577
rect 1170 12574 1176 12577
rect 712 12568 1176 12574
rect 1228 12574 1234 12577
rect 1686 12574 1692 12577
rect 1228 12568 1692 12574
rect 1744 12574 1750 12577
rect 2202 12574 2208 12577
rect 1744 12568 2208 12574
rect 2260 12574 2266 12577
rect 2718 12574 2724 12577
rect 2260 12568 2724 12574
rect 2776 12574 2782 12577
rect 3234 12574 3240 12577
rect 2776 12568 3240 12574
rect 3292 12574 3298 12577
rect 3750 12574 3756 12577
rect 3292 12568 3756 12574
rect 3808 12574 3814 12577
rect 4266 12574 4272 12577
rect 3808 12568 4272 12574
rect 4324 12574 4330 12577
rect 4782 12574 4788 12577
rect 4324 12568 4788 12574
rect 4840 12574 4846 12577
rect 5298 12574 5304 12577
rect 4840 12568 5304 12574
rect 5356 12574 5362 12577
rect 5814 12574 5820 12577
rect 5356 12568 5820 12574
rect 5872 12574 5878 12577
rect 6330 12574 6336 12577
rect 5872 12568 6336 12574
rect 6388 12574 6394 12577
rect 6846 12574 6852 12577
rect 6388 12568 6852 12574
rect 6904 12574 6910 12577
rect 7362 12574 7368 12577
rect 6904 12568 7368 12574
rect 7420 12574 7426 12577
rect 7878 12574 7884 12577
rect 7420 12568 7884 12574
rect 7936 12574 7942 12577
rect 8394 12574 8400 12577
rect 7936 12568 8400 12574
rect 8452 12574 8458 12577
rect 8910 12574 8916 12577
rect 8452 12568 8916 12574
rect 8968 12574 8974 12577
rect 9426 12574 9432 12577
rect 8968 12568 9432 12574
rect 9484 12574 9490 12577
rect 9942 12574 9948 12577
rect 9484 12568 9948 12574
rect 10000 12574 10006 12577
rect 10458 12574 10464 12577
rect 10000 12568 10464 12574
rect 10516 12574 10522 12577
rect 10974 12574 10980 12577
rect 10516 12568 10980 12574
rect 11032 12574 11038 12577
rect 11490 12574 11496 12577
rect 11032 12568 11496 12574
rect 11548 12574 11554 12577
rect 12006 12574 12012 12577
rect 11548 12568 12012 12574
rect 12064 12574 12070 12577
rect 12522 12574 12528 12577
rect 12064 12568 12528 12574
rect 12580 12574 12586 12577
rect 13038 12574 13044 12577
rect 12580 12568 13044 12574
rect 13096 12574 13102 12577
rect 13554 12574 13560 12577
rect 13096 12568 13560 12574
rect 13612 12574 13618 12577
rect 14070 12574 14076 12577
rect 13612 12568 14076 12574
rect 14128 12574 14134 12577
rect 14586 12574 14592 12577
rect 14128 12568 14592 12574
rect 14644 12574 14650 12577
rect 15102 12574 15108 12577
rect 14644 12568 15108 12574
rect 15160 12574 15166 12577
rect 15618 12574 15624 12577
rect 15160 12568 15624 12574
rect 15676 12574 15682 12577
rect 16134 12574 16140 12577
rect 15676 12568 16140 12574
rect 16192 12574 16198 12577
rect 16650 12574 16656 12577
rect 16192 12568 16656 12574
rect 16708 12574 16714 12577
rect 17166 12574 17172 12577
rect 16708 12568 17172 12574
rect 17224 12574 17230 12577
rect 17682 12574 17688 12577
rect 17224 12568 17688 12574
rect 17740 12574 17746 12577
rect 17740 12568 18129 12574
rect 271 12534 377 12568
rect 18023 12534 18129 12568
rect 271 12528 660 12534
rect 271 12468 317 12528
rect 654 12525 660 12528
rect 712 12528 1176 12534
rect 712 12525 718 12528
rect 1170 12525 1176 12528
rect 1228 12528 1692 12534
rect 1228 12525 1234 12528
rect 1686 12525 1692 12528
rect 1744 12528 2208 12534
rect 1744 12525 1750 12528
rect 2202 12525 2208 12528
rect 2260 12528 2724 12534
rect 2260 12525 2266 12528
rect 2718 12525 2724 12528
rect 2776 12528 3240 12534
rect 2776 12525 2782 12528
rect 3234 12525 3240 12528
rect 3292 12528 3756 12534
rect 3292 12525 3298 12528
rect 3750 12525 3756 12528
rect 3808 12528 4272 12534
rect 3808 12525 3814 12528
rect 4266 12525 4272 12528
rect 4324 12528 4788 12534
rect 4324 12525 4330 12528
rect 4782 12525 4788 12528
rect 4840 12528 5304 12534
rect 4840 12525 4846 12528
rect 5298 12525 5304 12528
rect 5356 12528 5820 12534
rect 5356 12525 5362 12528
rect 5814 12525 5820 12528
rect 5872 12528 6336 12534
rect 5872 12525 5878 12528
rect 6330 12525 6336 12528
rect 6388 12528 6852 12534
rect 6388 12525 6394 12528
rect 6846 12525 6852 12528
rect 6904 12528 7368 12534
rect 6904 12525 6910 12528
rect 7362 12525 7368 12528
rect 7420 12528 7884 12534
rect 7420 12525 7426 12528
rect 7878 12525 7884 12528
rect 7936 12528 8400 12534
rect 7936 12525 7942 12528
rect 8394 12525 8400 12528
rect 8452 12528 8916 12534
rect 8452 12525 8458 12528
rect 8910 12525 8916 12528
rect 8968 12528 9432 12534
rect 8968 12525 8974 12528
rect 9426 12525 9432 12528
rect 9484 12528 9948 12534
rect 9484 12525 9490 12528
rect 9942 12525 9948 12528
rect 10000 12528 10464 12534
rect 10000 12525 10006 12528
rect 10458 12525 10464 12528
rect 10516 12528 10980 12534
rect 10516 12525 10522 12528
rect 10974 12525 10980 12528
rect 11032 12528 11496 12534
rect 11032 12525 11038 12528
rect 11490 12525 11496 12528
rect 11548 12528 12012 12534
rect 11548 12525 11554 12528
rect 12006 12525 12012 12528
rect 12064 12528 12528 12534
rect 12064 12525 12070 12528
rect 12522 12525 12528 12528
rect 12580 12528 13044 12534
rect 12580 12525 12586 12528
rect 13038 12525 13044 12528
rect 13096 12528 13560 12534
rect 13096 12525 13102 12528
rect 13554 12525 13560 12528
rect 13612 12528 14076 12534
rect 13612 12525 13618 12528
rect 14070 12525 14076 12528
rect 14128 12528 14592 12534
rect 14128 12525 14134 12528
rect 14586 12525 14592 12528
rect 14644 12528 15108 12534
rect 14644 12525 14650 12528
rect 15102 12525 15108 12528
rect 15160 12528 15624 12534
rect 15160 12525 15166 12528
rect 15618 12525 15624 12528
rect 15676 12528 16140 12534
rect 15676 12525 15682 12528
rect 16134 12525 16140 12528
rect 16192 12528 16656 12534
rect 16192 12525 16198 12528
rect 16650 12525 16656 12528
rect 16708 12528 17172 12534
rect 16708 12525 16714 12528
rect 17166 12525 17172 12528
rect 17224 12528 17688 12534
rect 17224 12525 17230 12528
rect 17682 12525 17688 12528
rect 17740 12528 18129 12534
rect 17740 12525 17746 12528
rect 271 10730 277 12468
rect 311 10730 317 12468
rect 18083 12468 18129 12528
rect 402 12390 17998 12436
rect 402 12343 454 12390
rect 402 10808 454 10855
rect 660 12343 712 12349
rect 660 10849 712 10855
rect 918 12343 970 12349
rect 918 10849 970 10855
rect 1176 12343 1228 12349
rect 1176 10849 1228 10855
rect 1434 12343 1486 12349
rect 1434 10849 1486 10855
rect 1692 12343 1744 12349
rect 1692 10849 1744 10855
rect 1950 12343 2002 12349
rect 1950 10849 2002 10855
rect 2208 12343 2260 12349
rect 2208 10849 2260 10855
rect 2466 12343 2518 12349
rect 2466 10849 2518 10855
rect 2724 12343 2776 12349
rect 2724 10849 2776 10855
rect 2982 12343 3034 12349
rect 2982 10849 3034 10855
rect 3240 12343 3292 12349
rect 3240 10849 3292 10855
rect 3498 12343 3550 12349
rect 3498 10849 3550 10855
rect 3756 12343 3808 12349
rect 3756 10849 3808 10855
rect 4014 12343 4066 12349
rect 4014 10849 4066 10855
rect 4272 12343 4324 12349
rect 4272 10849 4324 10855
rect 4530 12343 4582 12349
rect 4530 10849 4582 10855
rect 4788 12343 4840 12349
rect 4788 10849 4840 10855
rect 5046 12343 5098 12349
rect 5046 10849 5098 10855
rect 5304 12343 5356 12349
rect 5304 10849 5356 10855
rect 5562 12343 5614 12349
rect 5562 10849 5614 10855
rect 5820 12343 5872 12349
rect 5820 10849 5872 10855
rect 6078 12343 6130 12349
rect 6078 10849 6130 10855
rect 6336 12343 6388 12349
rect 6336 10849 6388 10855
rect 6594 12343 6646 12349
rect 6594 10849 6646 10855
rect 6852 12343 6904 12349
rect 6852 10849 6904 10855
rect 7110 12343 7162 12349
rect 7110 10849 7162 10855
rect 7368 12343 7420 12349
rect 7368 10849 7420 10855
rect 7626 12343 7678 12349
rect 7626 10849 7678 10855
rect 7884 12343 7936 12349
rect 7884 10849 7936 10855
rect 8142 12343 8194 12349
rect 8142 10849 8194 10855
rect 8400 12343 8452 12349
rect 8400 10849 8452 10855
rect 8658 12343 8710 12349
rect 8658 10849 8710 10855
rect 8916 12343 8968 12349
rect 8916 10849 8968 10855
rect 9174 12343 9226 12390
rect 9174 10808 9226 10855
rect 9432 12343 9484 12349
rect 9432 10849 9484 10855
rect 9690 12343 9742 12349
rect 9690 10849 9742 10855
rect 9948 12343 10000 12349
rect 9948 10849 10000 10855
rect 10206 12343 10258 12349
rect 10206 10849 10258 10855
rect 10464 12343 10516 12349
rect 10464 10849 10516 10855
rect 10722 12343 10774 12349
rect 10722 10849 10774 10855
rect 10980 12343 11032 12349
rect 10980 10849 11032 10855
rect 11238 12343 11290 12349
rect 11238 10849 11290 10855
rect 11496 12343 11548 12349
rect 11496 10849 11548 10855
rect 11754 12343 11806 12349
rect 11754 10849 11806 10855
rect 12012 12343 12064 12349
rect 12012 10849 12064 10855
rect 12270 12343 12322 12349
rect 12270 10849 12322 10855
rect 12528 12343 12580 12349
rect 12528 10849 12580 10855
rect 12786 12343 12838 12349
rect 12786 10849 12838 10855
rect 13044 12343 13096 12349
rect 13044 10849 13096 10855
rect 13302 12343 13354 12349
rect 13302 10849 13354 10855
rect 13560 12343 13612 12349
rect 13560 10849 13612 10855
rect 13818 12343 13870 12349
rect 13818 10849 13870 10855
rect 14076 12343 14128 12349
rect 14076 10849 14128 10855
rect 14334 12343 14386 12349
rect 14334 10849 14386 10855
rect 14592 12343 14644 12349
rect 14592 10849 14644 10855
rect 14850 12343 14902 12349
rect 14850 10849 14902 10855
rect 15108 12343 15160 12349
rect 15108 10849 15160 10855
rect 15366 12343 15418 12349
rect 15366 10849 15418 10855
rect 15624 12343 15676 12349
rect 15624 10849 15676 10855
rect 15882 12343 15934 12349
rect 15882 10849 15934 10855
rect 16140 12343 16192 12349
rect 16140 10849 16192 10855
rect 16398 12343 16450 12349
rect 16398 10849 16450 10855
rect 16656 12343 16708 12349
rect 16656 10849 16708 10855
rect 16914 12343 16966 12349
rect 16914 10849 16966 10855
rect 17172 12343 17224 12349
rect 17172 10849 17224 10855
rect 17430 12343 17482 12349
rect 17430 10849 17482 10855
rect 17688 12343 17740 12349
rect 17688 10849 17740 10855
rect 17946 12343 17998 12390
rect 17946 10808 17998 10855
rect 402 10762 17998 10808
rect 271 10670 317 10730
rect 18083 10730 18089 12468
rect 18123 10730 18129 12468
rect 654 10670 660 10673
rect 271 10664 660 10670
rect 712 10670 718 10673
rect 1170 10670 1176 10673
rect 712 10664 1176 10670
rect 1228 10670 1234 10673
rect 1686 10670 1692 10673
rect 1228 10664 1692 10670
rect 1744 10670 1750 10673
rect 2202 10670 2208 10673
rect 1744 10664 2208 10670
rect 2260 10670 2266 10673
rect 2718 10670 2724 10673
rect 2260 10664 2724 10670
rect 2776 10670 2782 10673
rect 3234 10670 3240 10673
rect 2776 10664 3240 10670
rect 3292 10670 3298 10673
rect 3750 10670 3756 10673
rect 3292 10664 3756 10670
rect 3808 10670 3814 10673
rect 4266 10670 4272 10673
rect 3808 10664 4272 10670
rect 4324 10670 4330 10673
rect 4782 10670 4788 10673
rect 4324 10664 4788 10670
rect 4840 10670 4846 10673
rect 5298 10670 5304 10673
rect 4840 10664 5304 10670
rect 5356 10670 5362 10673
rect 5814 10670 5820 10673
rect 5356 10664 5820 10670
rect 5872 10670 5878 10673
rect 6330 10670 6336 10673
rect 5872 10664 6336 10670
rect 6388 10670 6394 10673
rect 6846 10670 6852 10673
rect 6388 10664 6852 10670
rect 6904 10670 6910 10673
rect 7362 10670 7368 10673
rect 6904 10664 7368 10670
rect 7420 10670 7426 10673
rect 7878 10670 7884 10673
rect 7420 10664 7884 10670
rect 7936 10670 7942 10673
rect 8394 10670 8400 10673
rect 7936 10664 8400 10670
rect 8452 10670 8458 10673
rect 8910 10670 8916 10673
rect 8452 10664 8916 10670
rect 8968 10670 8974 10673
rect 9426 10670 9432 10673
rect 8968 10664 9432 10670
rect 9484 10670 9490 10673
rect 9942 10670 9948 10673
rect 9484 10664 9948 10670
rect 10000 10670 10006 10673
rect 10458 10670 10464 10673
rect 10000 10664 10464 10670
rect 10516 10670 10522 10673
rect 10974 10670 10980 10673
rect 10516 10664 10980 10670
rect 11032 10670 11038 10673
rect 11490 10670 11496 10673
rect 11032 10664 11496 10670
rect 11548 10670 11554 10673
rect 12006 10670 12012 10673
rect 11548 10664 12012 10670
rect 12064 10670 12070 10673
rect 12522 10670 12528 10673
rect 12064 10664 12528 10670
rect 12580 10670 12586 10673
rect 13038 10670 13044 10673
rect 12580 10664 13044 10670
rect 13096 10670 13102 10673
rect 13554 10670 13560 10673
rect 13096 10664 13560 10670
rect 13612 10670 13618 10673
rect 14070 10670 14076 10673
rect 13612 10664 14076 10670
rect 14128 10670 14134 10673
rect 14586 10670 14592 10673
rect 14128 10664 14592 10670
rect 14644 10670 14650 10673
rect 15102 10670 15108 10673
rect 14644 10664 15108 10670
rect 15160 10670 15166 10673
rect 15618 10670 15624 10673
rect 15160 10664 15624 10670
rect 15676 10670 15682 10673
rect 16134 10670 16140 10673
rect 15676 10664 16140 10670
rect 16192 10670 16198 10673
rect 16650 10670 16656 10673
rect 16192 10664 16656 10670
rect 16708 10670 16714 10673
rect 17166 10670 17172 10673
rect 16708 10664 17172 10670
rect 17224 10670 17230 10673
rect 17682 10670 17688 10673
rect 17224 10664 17688 10670
rect 17740 10670 17746 10673
rect 18083 10670 18129 10730
rect 17740 10664 18129 10670
rect 271 10630 377 10664
rect 18023 10630 18129 10664
rect 271 10624 660 10630
rect 654 10621 660 10624
rect 712 10624 1176 10630
rect 712 10621 718 10624
rect 1170 10621 1176 10624
rect 1228 10624 1692 10630
rect 1228 10621 1234 10624
rect 1686 10621 1692 10624
rect 1744 10624 2208 10630
rect 1744 10621 1750 10624
rect 2202 10621 2208 10624
rect 2260 10624 2724 10630
rect 2260 10621 2266 10624
rect 2718 10621 2724 10624
rect 2776 10624 3240 10630
rect 2776 10621 2782 10624
rect 3234 10621 3240 10624
rect 3292 10624 3756 10630
rect 3292 10621 3298 10624
rect 3750 10621 3756 10624
rect 3808 10624 4272 10630
rect 3808 10621 3814 10624
rect 4266 10621 4272 10624
rect 4324 10624 4788 10630
rect 4324 10621 4330 10624
rect 4782 10621 4788 10624
rect 4840 10624 5304 10630
rect 4840 10621 4846 10624
rect 5298 10621 5304 10624
rect 5356 10624 5820 10630
rect 5356 10621 5362 10624
rect 5814 10621 5820 10624
rect 5872 10624 6336 10630
rect 5872 10621 5878 10624
rect 6330 10621 6336 10624
rect 6388 10624 6852 10630
rect 6388 10621 6394 10624
rect 6846 10621 6852 10624
rect 6904 10624 7368 10630
rect 6904 10621 6910 10624
rect 7362 10621 7368 10624
rect 7420 10624 7884 10630
rect 7420 10621 7426 10624
rect 7878 10621 7884 10624
rect 7936 10624 8400 10630
rect 7936 10621 7942 10624
rect 8394 10621 8400 10624
rect 8452 10624 8916 10630
rect 8452 10621 8458 10624
rect 8910 10621 8916 10624
rect 8968 10624 9432 10630
rect 8968 10621 8974 10624
rect 9426 10621 9432 10624
rect 9484 10624 9948 10630
rect 9484 10621 9490 10624
rect 9942 10621 9948 10624
rect 10000 10624 10464 10630
rect 10000 10621 10006 10624
rect 10458 10621 10464 10624
rect 10516 10624 10980 10630
rect 10516 10621 10522 10624
rect 10974 10621 10980 10624
rect 11032 10624 11496 10630
rect 11032 10621 11038 10624
rect 11490 10621 11496 10624
rect 11548 10624 12012 10630
rect 11548 10621 11554 10624
rect 12006 10621 12012 10624
rect 12064 10624 12528 10630
rect 12064 10621 12070 10624
rect 12522 10621 12528 10624
rect 12580 10624 13044 10630
rect 12580 10621 12586 10624
rect 13038 10621 13044 10624
rect 13096 10624 13560 10630
rect 13096 10621 13102 10624
rect 13554 10621 13560 10624
rect 13612 10624 14076 10630
rect 13612 10621 13618 10624
rect 14070 10621 14076 10624
rect 14128 10624 14592 10630
rect 14128 10621 14134 10624
rect 14586 10621 14592 10624
rect 14644 10624 15108 10630
rect 14644 10621 14650 10624
rect 15102 10621 15108 10624
rect 15160 10624 15624 10630
rect 15160 10621 15166 10624
rect 15618 10621 15624 10624
rect 15676 10624 16140 10630
rect 15676 10621 15682 10624
rect 16134 10621 16140 10624
rect 16192 10624 16656 10630
rect 16192 10621 16198 10624
rect 16650 10621 16656 10624
rect 16708 10624 17172 10630
rect 16708 10621 16714 10624
rect 17166 10621 17172 10624
rect 17224 10624 17688 10630
rect 17224 10621 17230 10624
rect 17682 10621 17688 10624
rect 17740 10624 18129 10630
rect 17740 10621 17746 10624
<< via1 >>
rect 660 12568 712 12577
rect 1176 12568 1228 12577
rect 1692 12568 1744 12577
rect 2208 12568 2260 12577
rect 2724 12568 2776 12577
rect 3240 12568 3292 12577
rect 3756 12568 3808 12577
rect 4272 12568 4324 12577
rect 4788 12568 4840 12577
rect 5304 12568 5356 12577
rect 5820 12568 5872 12577
rect 6336 12568 6388 12577
rect 6852 12568 6904 12577
rect 7368 12568 7420 12577
rect 7884 12568 7936 12577
rect 8400 12568 8452 12577
rect 8916 12568 8968 12577
rect 9432 12568 9484 12577
rect 9948 12568 10000 12577
rect 10464 12568 10516 12577
rect 10980 12568 11032 12577
rect 11496 12568 11548 12577
rect 12012 12568 12064 12577
rect 12528 12568 12580 12577
rect 13044 12568 13096 12577
rect 13560 12568 13612 12577
rect 14076 12568 14128 12577
rect 14592 12568 14644 12577
rect 15108 12568 15160 12577
rect 15624 12568 15676 12577
rect 16140 12568 16192 12577
rect 16656 12568 16708 12577
rect 17172 12568 17224 12577
rect 17688 12568 17740 12577
rect 660 12534 712 12568
rect 1176 12534 1228 12568
rect 1692 12534 1744 12568
rect 2208 12534 2260 12568
rect 2724 12534 2776 12568
rect 3240 12534 3292 12568
rect 3756 12534 3808 12568
rect 4272 12534 4324 12568
rect 4788 12534 4840 12568
rect 5304 12534 5356 12568
rect 5820 12534 5872 12568
rect 6336 12534 6388 12568
rect 6852 12534 6904 12568
rect 7368 12534 7420 12568
rect 7884 12534 7936 12568
rect 8400 12534 8452 12568
rect 8916 12534 8968 12568
rect 9432 12534 9484 12568
rect 9948 12534 10000 12568
rect 10464 12534 10516 12568
rect 10980 12534 11032 12568
rect 11496 12534 11548 12568
rect 12012 12534 12064 12568
rect 12528 12534 12580 12568
rect 13044 12534 13096 12568
rect 13560 12534 13612 12568
rect 14076 12534 14128 12568
rect 14592 12534 14644 12568
rect 15108 12534 15160 12568
rect 15624 12534 15676 12568
rect 16140 12534 16192 12568
rect 16656 12534 16708 12568
rect 17172 12534 17224 12568
rect 17688 12534 17740 12568
rect 660 12525 712 12534
rect 1176 12525 1228 12534
rect 1692 12525 1744 12534
rect 2208 12525 2260 12534
rect 2724 12525 2776 12534
rect 3240 12525 3292 12534
rect 3756 12525 3808 12534
rect 4272 12525 4324 12534
rect 4788 12525 4840 12534
rect 5304 12525 5356 12534
rect 5820 12525 5872 12534
rect 6336 12525 6388 12534
rect 6852 12525 6904 12534
rect 7368 12525 7420 12534
rect 7884 12525 7936 12534
rect 8400 12525 8452 12534
rect 8916 12525 8968 12534
rect 9432 12525 9484 12534
rect 9948 12525 10000 12534
rect 10464 12525 10516 12534
rect 10980 12525 11032 12534
rect 11496 12525 11548 12534
rect 12012 12525 12064 12534
rect 12528 12525 12580 12534
rect 13044 12525 13096 12534
rect 13560 12525 13612 12534
rect 14076 12525 14128 12534
rect 14592 12525 14644 12534
rect 15108 12525 15160 12534
rect 15624 12525 15676 12534
rect 16140 12525 16192 12534
rect 16656 12525 16708 12534
rect 17172 12525 17224 12534
rect 17688 12525 17740 12534
rect 402 10855 454 12343
rect 660 10855 712 12343
rect 918 10855 970 12343
rect 1176 10855 1228 12343
rect 1434 10855 1486 12343
rect 1692 10855 1744 12343
rect 1950 10855 2002 12343
rect 2208 10855 2260 12343
rect 2466 10855 2518 12343
rect 2724 10855 2776 12343
rect 2982 10855 3034 12343
rect 3240 10855 3292 12343
rect 3498 10855 3550 12343
rect 3756 10855 3808 12343
rect 4014 10855 4066 12343
rect 4272 10855 4324 12343
rect 4530 10855 4582 12343
rect 4788 10855 4840 12343
rect 5046 10855 5098 12343
rect 5304 10855 5356 12343
rect 5562 10855 5614 12343
rect 5820 10855 5872 12343
rect 6078 10855 6130 12343
rect 6336 10855 6388 12343
rect 6594 10855 6646 12343
rect 6852 10855 6904 12343
rect 7110 10855 7162 12343
rect 7368 10855 7420 12343
rect 7626 10855 7678 12343
rect 7884 10855 7936 12343
rect 8142 10855 8194 12343
rect 8400 10855 8452 12343
rect 8658 10855 8710 12343
rect 8916 10855 8968 12343
rect 9174 10855 9226 12343
rect 9432 10855 9484 12343
rect 9690 10855 9742 12343
rect 9948 10855 10000 12343
rect 10206 10855 10258 12343
rect 10464 10855 10516 12343
rect 10722 10855 10774 12343
rect 10980 10855 11032 12343
rect 11238 10855 11290 12343
rect 11496 10855 11548 12343
rect 11754 10855 11806 12343
rect 12012 10855 12064 12343
rect 12270 10855 12322 12343
rect 12528 10855 12580 12343
rect 12786 10855 12838 12343
rect 13044 10855 13096 12343
rect 13302 10855 13354 12343
rect 13560 10855 13612 12343
rect 13818 10855 13870 12343
rect 14076 10855 14128 12343
rect 14334 10855 14386 12343
rect 14592 10855 14644 12343
rect 14850 10855 14902 12343
rect 15108 10855 15160 12343
rect 15366 10855 15418 12343
rect 15624 10855 15676 12343
rect 15882 10855 15934 12343
rect 16140 10855 16192 12343
rect 16398 10855 16450 12343
rect 16656 10855 16708 12343
rect 16914 10855 16966 12343
rect 17172 10855 17224 12343
rect 17430 10855 17482 12343
rect 17688 10855 17740 12343
rect 17946 10855 17998 12343
rect 660 10664 712 10673
rect 1176 10664 1228 10673
rect 1692 10664 1744 10673
rect 2208 10664 2260 10673
rect 2724 10664 2776 10673
rect 3240 10664 3292 10673
rect 3756 10664 3808 10673
rect 4272 10664 4324 10673
rect 4788 10664 4840 10673
rect 5304 10664 5356 10673
rect 5820 10664 5872 10673
rect 6336 10664 6388 10673
rect 6852 10664 6904 10673
rect 7368 10664 7420 10673
rect 7884 10664 7936 10673
rect 8400 10664 8452 10673
rect 8916 10664 8968 10673
rect 9432 10664 9484 10673
rect 9948 10664 10000 10673
rect 10464 10664 10516 10673
rect 10980 10664 11032 10673
rect 11496 10664 11548 10673
rect 12012 10664 12064 10673
rect 12528 10664 12580 10673
rect 13044 10664 13096 10673
rect 13560 10664 13612 10673
rect 14076 10664 14128 10673
rect 14592 10664 14644 10673
rect 15108 10664 15160 10673
rect 15624 10664 15676 10673
rect 16140 10664 16192 10673
rect 16656 10664 16708 10673
rect 17172 10664 17224 10673
rect 17688 10664 17740 10673
rect 660 10630 712 10664
rect 1176 10630 1228 10664
rect 1692 10630 1744 10664
rect 2208 10630 2260 10664
rect 2724 10630 2776 10664
rect 3240 10630 3292 10664
rect 3756 10630 3808 10664
rect 4272 10630 4324 10664
rect 4788 10630 4840 10664
rect 5304 10630 5356 10664
rect 5820 10630 5872 10664
rect 6336 10630 6388 10664
rect 6852 10630 6904 10664
rect 7368 10630 7420 10664
rect 7884 10630 7936 10664
rect 8400 10630 8452 10664
rect 8916 10630 8968 10664
rect 9432 10630 9484 10664
rect 9948 10630 10000 10664
rect 10464 10630 10516 10664
rect 10980 10630 11032 10664
rect 11496 10630 11548 10664
rect 12012 10630 12064 10664
rect 12528 10630 12580 10664
rect 13044 10630 13096 10664
rect 13560 10630 13612 10664
rect 14076 10630 14128 10664
rect 14592 10630 14644 10664
rect 15108 10630 15160 10664
rect 15624 10630 15676 10664
rect 16140 10630 16192 10664
rect 16656 10630 16708 10664
rect 17172 10630 17224 10664
rect 17688 10630 17740 10664
rect 660 10621 712 10630
rect 1176 10621 1228 10630
rect 1692 10621 1744 10630
rect 2208 10621 2260 10630
rect 2724 10621 2776 10630
rect 3240 10621 3292 10630
rect 3756 10621 3808 10630
rect 4272 10621 4324 10630
rect 4788 10621 4840 10630
rect 5304 10621 5356 10630
rect 5820 10621 5872 10630
rect 6336 10621 6388 10630
rect 6852 10621 6904 10630
rect 7368 10621 7420 10630
rect 7884 10621 7936 10630
rect 8400 10621 8452 10630
rect 8916 10621 8968 10630
rect 9432 10621 9484 10630
rect 9948 10621 10000 10630
rect 10464 10621 10516 10630
rect 10980 10621 11032 10630
rect 11496 10621 11548 10630
rect 12012 10621 12064 10630
rect 12528 10621 12580 10630
rect 13044 10621 13096 10630
rect 13560 10621 13612 10630
rect 14076 10621 14128 10630
rect 14592 10621 14644 10630
rect 15108 10621 15160 10630
rect 15624 10621 15676 10630
rect 16140 10621 16192 10630
rect 16656 10621 16708 10630
rect 17172 10621 17224 10630
rect 17688 10621 17740 10630
<< metal2 >>
rect 351 12879 505 12884
rect 351 12739 360 12879
rect 496 12739 505 12879
rect 351 12734 505 12739
rect 402 12343 454 12734
rect 654 12525 660 12577
rect 712 12525 718 12577
rect 660 12343 712 12525
rect 618 11779 660 11788
rect 918 12343 970 12884
rect 1170 12525 1176 12577
rect 1228 12525 1234 12577
rect 712 11779 754 11788
rect 618 11410 660 11419
rect 402 10314 454 10855
rect 712 11410 754 11419
rect 660 10673 712 10855
rect 1176 12343 1228 12525
rect 1134 11779 1176 11788
rect 1434 12343 1486 12884
rect 1686 12525 1692 12577
rect 1744 12525 1750 12577
rect 1228 11779 1270 11788
rect 1134 11410 1176 11419
rect 654 10621 660 10673
rect 712 10621 718 10673
rect 918 10464 970 10855
rect 1228 11410 1270 11419
rect 1176 10673 1228 10855
rect 1692 12343 1744 12525
rect 1950 12444 2002 12884
rect 2202 12525 2208 12577
rect 2260 12525 2266 12577
rect 1650 11779 1692 11788
rect 1899 12439 2053 12444
rect 1899 12299 1908 12439
rect 2044 12299 2053 12439
rect 1899 12294 1950 12299
rect 1744 11779 1786 11788
rect 1650 11410 1692 11419
rect 1434 10684 1486 10855
rect 1744 11410 1786 11419
rect 1383 10679 1537 10684
rect 1170 10621 1176 10673
rect 1228 10621 1234 10673
rect 1383 10539 1392 10679
rect 1528 10539 1537 10679
rect 1692 10673 1744 10855
rect 2002 12294 2053 12299
rect 2208 12343 2260 12525
rect 2166 11779 2208 11788
rect 2466 12343 2518 12884
rect 2982 12664 3034 12884
rect 3498 12664 3550 12884
rect 2931 12659 3085 12664
rect 2718 12525 2724 12577
rect 2776 12525 2782 12577
rect 2260 11779 2302 11788
rect 2166 11410 2208 11419
rect 1686 10621 1692 10673
rect 1744 10621 1750 10673
rect 1383 10534 1537 10539
rect 867 10459 1021 10464
rect 867 10319 876 10459
rect 1012 10319 1021 10459
rect 867 10314 1021 10319
rect 1434 10314 1486 10534
rect 1950 10314 2002 10855
rect 2260 11410 2302 11419
rect 2208 10673 2260 10855
rect 2415 10899 2466 10904
rect 2724 12343 2776 12525
rect 2931 12519 2940 12659
rect 3076 12519 3085 12659
rect 3447 12659 3601 12664
rect 3234 12525 3240 12577
rect 3292 12525 3298 12577
rect 2931 12514 3085 12519
rect 2682 11779 2724 11788
rect 2982 12343 3034 12514
rect 2776 11779 2818 11788
rect 2682 11410 2724 11419
rect 2518 10899 2569 10904
rect 2415 10759 2424 10899
rect 2560 10759 2569 10899
rect 2415 10754 2569 10759
rect 2776 11410 2818 11419
rect 2202 10621 2208 10673
rect 2260 10621 2266 10673
rect 2466 10314 2518 10754
rect 2724 10673 2776 10855
rect 3240 12343 3292 12525
rect 3447 12519 3456 12659
rect 3592 12519 3601 12659
rect 3750 12525 3756 12577
rect 3808 12525 3814 12577
rect 3447 12514 3601 12519
rect 3198 11779 3240 11788
rect 3498 12343 3550 12514
rect 3292 11779 3334 11788
rect 3198 11410 3240 11419
rect 2718 10621 2724 10673
rect 2776 10621 2782 10673
rect 2982 10314 3034 10855
rect 3292 11410 3334 11419
rect 3240 10673 3292 10855
rect 3756 12343 3808 12525
rect 3714 11779 3756 11788
rect 4014 12343 4066 12884
rect 4266 12525 4272 12577
rect 4324 12525 4330 12577
rect 3808 11779 3850 11788
rect 3714 11410 3756 11419
rect 3234 10621 3240 10673
rect 3292 10621 3298 10673
rect 3498 10314 3550 10855
rect 3808 11410 3850 11419
rect 3963 11339 4014 11344
rect 4272 12343 4324 12525
rect 4230 11779 4272 11788
rect 4530 12343 4582 12884
rect 4782 12525 4788 12577
rect 4840 12525 4846 12577
rect 4479 11999 4530 12004
rect 4788 12343 4840 12525
rect 4582 11999 4633 12004
rect 4479 11859 4488 11999
rect 4624 11859 4633 11999
rect 4479 11854 4530 11859
rect 4324 11779 4366 11788
rect 4230 11410 4272 11419
rect 4066 11339 4117 11344
rect 3963 11199 3972 11339
rect 4108 11199 4117 11339
rect 3963 11194 4014 11199
rect 3756 10673 3808 10855
rect 4066 11194 4117 11199
rect 3750 10621 3756 10673
rect 3808 10621 3814 10673
rect 4014 10314 4066 10855
rect 4324 11410 4366 11419
rect 4272 10673 4324 10855
rect 4582 11854 4633 11859
rect 4746 11779 4788 11788
rect 5046 12343 5098 12884
rect 5298 12525 5304 12577
rect 5356 12525 5362 12577
rect 4840 11779 4882 11788
rect 4746 11410 4788 11419
rect 4266 10621 4272 10673
rect 4324 10621 4330 10673
rect 4530 10314 4582 10855
rect 4840 11410 4882 11419
rect 4788 10673 4840 10855
rect 5304 12343 5356 12525
rect 5262 11779 5304 11788
rect 5562 12343 5614 12884
rect 5814 12525 5820 12577
rect 5872 12525 5878 12577
rect 5356 11779 5398 11788
rect 5262 11410 5304 11419
rect 4782 10621 4788 10673
rect 4840 10621 4846 10673
rect 5046 10464 5098 10855
rect 5356 11410 5398 11419
rect 5304 10673 5356 10855
rect 5820 12343 5872 12525
rect 5778 11779 5820 11788
rect 6078 12343 6130 12884
rect 6330 12525 6336 12577
rect 6388 12525 6394 12577
rect 6027 12219 6078 12224
rect 6336 12343 6388 12525
rect 6130 12219 6181 12224
rect 6027 12079 6036 12219
rect 6172 12079 6181 12219
rect 6027 12074 6078 12079
rect 5872 11779 5914 11788
rect 5778 11410 5820 11419
rect 5562 10684 5614 10855
rect 5872 11410 5914 11419
rect 5511 10679 5665 10684
rect 5298 10621 5304 10673
rect 5356 10621 5362 10673
rect 5511 10539 5520 10679
rect 5656 10539 5665 10679
rect 5820 10673 5872 10855
rect 6130 12074 6181 12079
rect 6294 11779 6336 11788
rect 6594 12343 6646 12884
rect 7110 12664 7162 12884
rect 7626 12664 7678 12884
rect 7059 12659 7213 12664
rect 6846 12525 6852 12577
rect 6904 12525 6910 12577
rect 6388 11779 6430 11788
rect 6294 11410 6336 11419
rect 5814 10621 5820 10673
rect 5872 10621 5878 10673
rect 5511 10534 5665 10539
rect 4995 10459 5149 10464
rect 4995 10319 5004 10459
rect 5140 10319 5149 10459
rect 4995 10314 5149 10319
rect 5562 10314 5614 10534
rect 6078 10314 6130 10855
rect 6388 11410 6430 11419
rect 6543 11119 6594 11124
rect 6852 12343 6904 12525
rect 7059 12519 7068 12659
rect 7204 12519 7213 12659
rect 7575 12659 7729 12664
rect 7362 12525 7368 12577
rect 7420 12525 7426 12577
rect 7059 12514 7213 12519
rect 6810 11779 6852 11788
rect 7110 12343 7162 12514
rect 6904 11779 6946 11788
rect 6810 11410 6852 11419
rect 6646 11119 6697 11124
rect 6543 10979 6552 11119
rect 6688 10979 6697 11119
rect 6543 10974 6594 10979
rect 6336 10673 6388 10855
rect 6646 10974 6697 10979
rect 6330 10621 6336 10673
rect 6388 10621 6394 10673
rect 6594 10314 6646 10855
rect 6904 11410 6946 11419
rect 6852 10673 6904 10855
rect 7368 12343 7420 12525
rect 7575 12519 7584 12659
rect 7720 12519 7729 12659
rect 7878 12525 7884 12577
rect 7936 12525 7942 12577
rect 7575 12514 7729 12519
rect 7326 11779 7368 11788
rect 7626 12343 7678 12514
rect 7420 11779 7462 11788
rect 7326 11410 7368 11419
rect 6846 10621 6852 10673
rect 6904 10621 6910 10673
rect 7110 10314 7162 10855
rect 7420 11410 7462 11419
rect 7368 10673 7420 10855
rect 7884 12343 7936 12525
rect 7842 11779 7884 11788
rect 8142 12343 8194 12884
rect 8394 12525 8400 12577
rect 8452 12525 8458 12577
rect 7936 11779 7978 11788
rect 7842 11410 7884 11419
rect 7362 10621 7368 10673
rect 7420 10621 7426 10673
rect 7626 10314 7678 10855
rect 7936 11410 7978 11419
rect 8091 11339 8142 11344
rect 8400 12343 8452 12525
rect 8358 11779 8400 11788
rect 8658 12343 8710 12884
rect 9123 12879 9277 12884
rect 9123 12739 9132 12879
rect 9268 12739 9277 12879
rect 9123 12734 9277 12739
rect 8910 12525 8916 12577
rect 8968 12525 8974 12577
rect 8607 11999 8658 12004
rect 8916 12343 8968 12525
rect 8710 11999 8761 12004
rect 8607 11859 8616 11999
rect 8752 11859 8761 11999
rect 8607 11854 8658 11859
rect 8452 11779 8494 11788
rect 8358 11410 8400 11419
rect 8194 11339 8245 11344
rect 8091 11199 8100 11339
rect 8236 11199 8245 11339
rect 8091 11194 8142 11199
rect 7884 10673 7936 10855
rect 8194 11194 8245 11199
rect 7878 10621 7884 10673
rect 7936 10621 7942 10673
rect 8142 10314 8194 10855
rect 8452 11410 8494 11419
rect 8400 10673 8452 10855
rect 8710 11854 8761 11859
rect 8874 11779 8916 11788
rect 9174 12343 9226 12734
rect 9426 12525 9432 12577
rect 9484 12525 9490 12577
rect 8968 11779 9010 11788
rect 8874 11410 8916 11419
rect 8394 10621 8400 10673
rect 8452 10621 8458 10673
rect 8658 10314 8710 10855
rect 8968 11410 9010 11419
rect 8916 10673 8968 10855
rect 9432 12343 9484 12525
rect 9390 11779 9432 11788
rect 9690 12343 9742 12884
rect 9942 12525 9948 12577
rect 10000 12525 10006 12577
rect 9639 11999 9690 12004
rect 9948 12343 10000 12525
rect 9742 11999 9793 12004
rect 9639 11859 9648 11999
rect 9784 11859 9793 11999
rect 9639 11854 9690 11859
rect 9484 11779 9526 11788
rect 9390 11410 9432 11419
rect 8910 10621 8916 10673
rect 8968 10621 8974 10673
rect 9174 10314 9226 10855
rect 9484 11410 9526 11419
rect 9432 10673 9484 10855
rect 9742 11854 9793 11859
rect 9906 11779 9948 11788
rect 10206 12343 10258 12884
rect 10722 12664 10774 12884
rect 11238 12664 11290 12884
rect 10671 12659 10825 12664
rect 10458 12525 10464 12577
rect 10516 12525 10522 12577
rect 10000 11779 10042 11788
rect 9906 11410 9948 11419
rect 9426 10621 9432 10673
rect 9484 10621 9490 10673
rect 9690 10314 9742 10855
rect 10000 11410 10042 11419
rect 10155 11339 10206 11344
rect 10464 12343 10516 12525
rect 10671 12519 10680 12659
rect 10816 12519 10825 12659
rect 11187 12659 11341 12664
rect 10974 12525 10980 12577
rect 11032 12525 11038 12577
rect 10671 12514 10825 12519
rect 10422 11779 10464 11788
rect 10722 12343 10774 12514
rect 10516 11779 10558 11788
rect 10422 11410 10464 11419
rect 10258 11339 10309 11344
rect 10155 11199 10164 11339
rect 10300 11199 10309 11339
rect 10155 11194 10206 11199
rect 9948 10673 10000 10855
rect 10258 11194 10309 11199
rect 9942 10621 9948 10673
rect 10000 10621 10006 10673
rect 10206 10314 10258 10855
rect 10516 11410 10558 11419
rect 10464 10673 10516 10855
rect 10980 12343 11032 12525
rect 11187 12519 11196 12659
rect 11332 12519 11341 12659
rect 11490 12525 11496 12577
rect 11548 12525 11554 12577
rect 11187 12514 11341 12519
rect 10938 11779 10980 11788
rect 11238 12343 11290 12514
rect 11032 11779 11074 11788
rect 10938 11410 10980 11419
rect 10458 10621 10464 10673
rect 10516 10621 10522 10673
rect 10722 10314 10774 10855
rect 11032 11410 11074 11419
rect 10980 10673 11032 10855
rect 11496 12343 11548 12525
rect 11454 11779 11496 11788
rect 11754 12343 11806 12884
rect 12006 12525 12012 12577
rect 12064 12525 12070 12577
rect 11548 11779 11590 11788
rect 11454 11410 11496 11419
rect 10974 10621 10980 10673
rect 11032 10621 11038 10673
rect 11238 10314 11290 10855
rect 11548 11410 11590 11419
rect 11703 11119 11754 11124
rect 12012 12343 12064 12525
rect 11970 11779 12012 11788
rect 12270 12343 12322 12884
rect 12522 12525 12528 12577
rect 12580 12525 12586 12577
rect 12219 12219 12270 12224
rect 12528 12343 12580 12525
rect 12322 12219 12373 12224
rect 12219 12079 12228 12219
rect 12364 12079 12373 12219
rect 12219 12074 12270 12079
rect 12064 11779 12106 11788
rect 11970 11410 12012 11419
rect 11806 11119 11857 11124
rect 11703 10979 11712 11119
rect 11848 10979 11857 11119
rect 11703 10974 11754 10979
rect 11496 10673 11548 10855
rect 11806 10974 11857 10979
rect 11490 10621 11496 10673
rect 11548 10621 11554 10673
rect 11754 10314 11806 10855
rect 12064 11410 12106 11419
rect 12012 10673 12064 10855
rect 12322 12074 12373 12079
rect 12486 11779 12528 11788
rect 12786 12343 12838 12884
rect 13038 12525 13044 12577
rect 13096 12525 13102 12577
rect 12580 11779 12622 11788
rect 12486 11410 12528 11419
rect 12006 10621 12012 10673
rect 12064 10621 12070 10673
rect 12270 10314 12322 10855
rect 12580 11410 12622 11419
rect 12528 10673 12580 10855
rect 13044 12343 13096 12525
rect 13002 11779 13044 11788
rect 13302 12343 13354 12884
rect 13554 12525 13560 12577
rect 13612 12525 13618 12577
rect 13096 11779 13138 11788
rect 13002 11410 13044 11419
rect 12786 10684 12838 10855
rect 13096 11410 13138 11419
rect 12735 10679 12889 10684
rect 12522 10621 12528 10673
rect 12580 10621 12586 10673
rect 12735 10539 12744 10679
rect 12880 10539 12889 10679
rect 13044 10673 13096 10855
rect 13560 12343 13612 12525
rect 13518 11779 13560 11788
rect 13818 12343 13870 12884
rect 14070 12525 14076 12577
rect 14128 12525 14134 12577
rect 13767 11999 13818 12004
rect 14076 12343 14128 12525
rect 13870 11999 13921 12004
rect 13767 11859 13776 11999
rect 13912 11859 13921 11999
rect 13767 11854 13818 11859
rect 13612 11779 13654 11788
rect 13518 11410 13560 11419
rect 13038 10621 13044 10673
rect 13096 10621 13102 10673
rect 12735 10534 12889 10539
rect 12786 10314 12838 10534
rect 13302 10464 13354 10855
rect 13612 11410 13654 11419
rect 13560 10673 13612 10855
rect 13870 11854 13921 11859
rect 14034 11779 14076 11788
rect 14334 12343 14386 12884
rect 14850 12664 14902 12884
rect 15366 12664 15418 12884
rect 14799 12659 14953 12664
rect 14586 12525 14592 12577
rect 14644 12525 14650 12577
rect 14128 11779 14170 11788
rect 14034 11410 14076 11419
rect 13554 10621 13560 10673
rect 13612 10621 13618 10673
rect 13251 10459 13405 10464
rect 13251 10319 13260 10459
rect 13396 10319 13405 10459
rect 13251 10314 13405 10319
rect 13818 10314 13870 10855
rect 14128 11410 14170 11419
rect 14283 11339 14334 11344
rect 14592 12343 14644 12525
rect 14799 12519 14808 12659
rect 14944 12519 14953 12659
rect 15315 12659 15469 12664
rect 15102 12525 15108 12577
rect 15160 12525 15166 12577
rect 14799 12514 14953 12519
rect 14550 11779 14592 11788
rect 14850 12343 14902 12514
rect 14644 11779 14686 11788
rect 14550 11410 14592 11419
rect 14386 11339 14437 11344
rect 14283 11199 14292 11339
rect 14428 11199 14437 11339
rect 14283 11194 14334 11199
rect 14076 10673 14128 10855
rect 14386 11194 14437 11199
rect 14070 10621 14076 10673
rect 14128 10621 14134 10673
rect 14334 10314 14386 10855
rect 14644 11410 14686 11419
rect 14592 10673 14644 10855
rect 15108 12343 15160 12525
rect 15315 12519 15324 12659
rect 15460 12519 15469 12659
rect 15618 12525 15624 12577
rect 15676 12525 15682 12577
rect 15315 12514 15469 12519
rect 15066 11779 15108 11788
rect 15366 12343 15418 12514
rect 15160 11779 15202 11788
rect 15066 11410 15108 11419
rect 14586 10621 14592 10673
rect 14644 10621 14650 10673
rect 14850 10314 14902 10855
rect 15160 11410 15202 11419
rect 15108 10673 15160 10855
rect 15624 12343 15676 12525
rect 15582 11779 15624 11788
rect 15882 12343 15934 12884
rect 16134 12525 16140 12577
rect 16192 12525 16198 12577
rect 15676 11779 15718 11788
rect 15582 11410 15624 11419
rect 15102 10621 15108 10673
rect 15160 10621 15166 10673
rect 15366 10314 15418 10855
rect 15676 11410 15718 11419
rect 15624 10673 15676 10855
rect 15831 10899 15882 10904
rect 16140 12343 16192 12525
rect 16398 12444 16450 12884
rect 16650 12525 16656 12577
rect 16708 12525 16714 12577
rect 16098 11779 16140 11788
rect 16347 12439 16501 12444
rect 16347 12299 16356 12439
rect 16492 12299 16501 12439
rect 16347 12294 16398 12299
rect 16192 11779 16234 11788
rect 16098 11410 16140 11419
rect 15934 10899 15985 10904
rect 15831 10759 15840 10899
rect 15976 10759 15985 10899
rect 15831 10754 15985 10759
rect 16192 11410 16234 11419
rect 15618 10621 15624 10673
rect 15676 10621 15682 10673
rect 15882 10314 15934 10754
rect 16140 10673 16192 10855
rect 16450 12294 16501 12299
rect 16656 12343 16708 12525
rect 16614 11779 16656 11788
rect 16914 12343 16966 12884
rect 17166 12525 17172 12577
rect 17224 12525 17230 12577
rect 16708 11779 16750 11788
rect 16614 11410 16656 11419
rect 16134 10621 16140 10673
rect 16192 10621 16198 10673
rect 16398 10314 16450 10855
rect 16708 11410 16750 11419
rect 16656 10673 16708 10855
rect 17172 12343 17224 12525
rect 17130 11779 17172 11788
rect 17430 12343 17482 12884
rect 17895 12879 18049 12884
rect 17895 12739 17904 12879
rect 18040 12739 18049 12879
rect 17895 12734 18049 12739
rect 17682 12525 17688 12577
rect 17740 12525 17746 12577
rect 17224 11779 17266 11788
rect 17130 11410 17172 11419
rect 16914 10684 16966 10855
rect 17224 11410 17266 11419
rect 16863 10679 17017 10684
rect 16650 10621 16656 10673
rect 16708 10621 16714 10673
rect 16863 10539 16872 10679
rect 17008 10539 17017 10679
rect 17172 10673 17224 10855
rect 17688 12343 17740 12525
rect 17646 11779 17688 11788
rect 17946 12343 17998 12734
rect 17740 11779 17782 11788
rect 17646 11410 17688 11419
rect 17166 10621 17172 10673
rect 17224 10621 17230 10673
rect 16863 10534 17017 10539
rect 16914 10314 16966 10534
rect 17430 10464 17482 10855
rect 17740 11410 17782 11419
rect 17688 10673 17740 10855
rect 17682 10621 17688 10673
rect 17740 10621 17746 10673
rect 17379 10459 17533 10464
rect 17379 10319 17388 10459
rect 17524 10319 17533 10459
rect 17379 10314 17533 10319
rect 17946 10314 17998 10855
<< via2 >>
rect 360 12739 496 12879
rect 618 11419 660 11779
rect 660 11419 712 11779
rect 712 11419 754 11779
rect 1134 11419 1176 11779
rect 1176 11419 1228 11779
rect 1228 11419 1270 11779
rect 1908 12343 2044 12439
rect 1908 12299 1950 12343
rect 1950 12299 2002 12343
rect 2002 12299 2044 12343
rect 1650 11419 1692 11779
rect 1692 11419 1744 11779
rect 1744 11419 1786 11779
rect 1392 10539 1528 10679
rect 2166 11419 2208 11779
rect 2208 11419 2260 11779
rect 2260 11419 2302 11779
rect 876 10319 1012 10459
rect 2940 12519 3076 12659
rect 2682 11419 2724 11779
rect 2724 11419 2776 11779
rect 2776 11419 2818 11779
rect 2424 10855 2466 10899
rect 2466 10855 2518 10899
rect 2518 10855 2560 10899
rect 2424 10759 2560 10855
rect 3456 12519 3592 12659
rect 3198 11419 3240 11779
rect 3240 11419 3292 11779
rect 3292 11419 3334 11779
rect 3714 11419 3756 11779
rect 3756 11419 3808 11779
rect 3808 11419 3850 11779
rect 4488 11859 4530 11999
rect 4530 11859 4582 11999
rect 4582 11859 4624 11999
rect 4230 11419 4272 11779
rect 4272 11419 4324 11779
rect 4324 11419 4366 11779
rect 3972 11199 4014 11339
rect 4014 11199 4066 11339
rect 4066 11199 4108 11339
rect 4746 11419 4788 11779
rect 4788 11419 4840 11779
rect 4840 11419 4882 11779
rect 5262 11419 5304 11779
rect 5304 11419 5356 11779
rect 5356 11419 5398 11779
rect 6036 12079 6078 12219
rect 6078 12079 6130 12219
rect 6130 12079 6172 12219
rect 5778 11419 5820 11779
rect 5820 11419 5872 11779
rect 5872 11419 5914 11779
rect 5520 10539 5656 10679
rect 6294 11419 6336 11779
rect 6336 11419 6388 11779
rect 6388 11419 6430 11779
rect 5004 10319 5140 10459
rect 7068 12519 7204 12659
rect 6810 11419 6852 11779
rect 6852 11419 6904 11779
rect 6904 11419 6946 11779
rect 6552 10979 6594 11119
rect 6594 10979 6646 11119
rect 6646 10979 6688 11119
rect 7584 12519 7720 12659
rect 7326 11419 7368 11779
rect 7368 11419 7420 11779
rect 7420 11419 7462 11779
rect 7842 11419 7884 11779
rect 7884 11419 7936 11779
rect 7936 11419 7978 11779
rect 9132 12739 9268 12879
rect 8616 11859 8658 11999
rect 8658 11859 8710 11999
rect 8710 11859 8752 11999
rect 8358 11419 8400 11779
rect 8400 11419 8452 11779
rect 8452 11419 8494 11779
rect 8100 11199 8142 11339
rect 8142 11199 8194 11339
rect 8194 11199 8236 11339
rect 8874 11419 8916 11779
rect 8916 11419 8968 11779
rect 8968 11419 9010 11779
rect 9648 11859 9690 11999
rect 9690 11859 9742 11999
rect 9742 11859 9784 11999
rect 9390 11419 9432 11779
rect 9432 11419 9484 11779
rect 9484 11419 9526 11779
rect 9906 11419 9948 11779
rect 9948 11419 10000 11779
rect 10000 11419 10042 11779
rect 10680 12519 10816 12659
rect 10422 11419 10464 11779
rect 10464 11419 10516 11779
rect 10516 11419 10558 11779
rect 10164 11199 10206 11339
rect 10206 11199 10258 11339
rect 10258 11199 10300 11339
rect 11196 12519 11332 12659
rect 10938 11419 10980 11779
rect 10980 11419 11032 11779
rect 11032 11419 11074 11779
rect 11454 11419 11496 11779
rect 11496 11419 11548 11779
rect 11548 11419 11590 11779
rect 12228 12079 12270 12219
rect 12270 12079 12322 12219
rect 12322 12079 12364 12219
rect 11970 11419 12012 11779
rect 12012 11419 12064 11779
rect 12064 11419 12106 11779
rect 11712 10979 11754 11119
rect 11754 10979 11806 11119
rect 11806 10979 11848 11119
rect 12486 11419 12528 11779
rect 12528 11419 12580 11779
rect 12580 11419 12622 11779
rect 13002 11419 13044 11779
rect 13044 11419 13096 11779
rect 13096 11419 13138 11779
rect 12744 10539 12880 10679
rect 13776 11859 13818 11999
rect 13818 11859 13870 11999
rect 13870 11859 13912 11999
rect 13518 11419 13560 11779
rect 13560 11419 13612 11779
rect 13612 11419 13654 11779
rect 14034 11419 14076 11779
rect 14076 11419 14128 11779
rect 14128 11419 14170 11779
rect 13260 10319 13396 10459
rect 14808 12519 14944 12659
rect 14550 11419 14592 11779
rect 14592 11419 14644 11779
rect 14644 11419 14686 11779
rect 14292 11199 14334 11339
rect 14334 11199 14386 11339
rect 14386 11199 14428 11339
rect 15324 12519 15460 12659
rect 15066 11419 15108 11779
rect 15108 11419 15160 11779
rect 15160 11419 15202 11779
rect 15582 11419 15624 11779
rect 15624 11419 15676 11779
rect 15676 11419 15718 11779
rect 16356 12343 16492 12439
rect 16356 12299 16398 12343
rect 16398 12299 16450 12343
rect 16450 12299 16492 12343
rect 16098 11419 16140 11779
rect 16140 11419 16192 11779
rect 16192 11419 16234 11779
rect 15840 10855 15882 10899
rect 15882 10855 15934 10899
rect 15934 10855 15976 10899
rect 15840 10759 15976 10855
rect 16614 11419 16656 11779
rect 16656 11419 16708 11779
rect 16708 11419 16750 11779
rect 17904 12739 18040 12879
rect 17130 11419 17172 11779
rect 17172 11419 17224 11779
rect 17224 11419 17266 11779
rect 16872 10539 17008 10679
rect 17646 11419 17688 11779
rect 17688 11419 17740 11779
rect 17740 11419 17782 11779
rect 17388 10319 17524 10459
<< metal3 >>
rect 20 12879 18380 12884
rect 20 12739 360 12879
rect 496 12739 9132 12879
rect 9268 12739 17904 12879
rect 18040 12739 18380 12879
rect 20 12734 18380 12739
rect 20 12663 18380 12664
rect 20 12659 13331 12663
rect 20 12519 2940 12659
rect 3076 12519 3456 12659
rect 3592 12519 7068 12659
rect 7204 12519 7584 12659
rect 7720 12519 10680 12659
rect 10816 12519 11196 12659
rect 11332 12519 13331 12659
rect 20 12515 13331 12519
rect 13629 12659 18380 12663
rect 13629 12519 14808 12659
rect 14944 12519 15324 12659
rect 15460 12519 18380 12659
rect 13629 12515 18380 12519
rect 20 12514 18380 12515
rect 20 12443 18380 12444
rect 20 12439 9051 12443
rect 20 12299 1908 12439
rect 2044 12299 9051 12439
rect 20 12295 9051 12299
rect 9349 12439 18380 12443
rect 9349 12299 16356 12439
rect 16492 12299 18380 12439
rect 9349 12295 18380 12299
rect 20 12294 18380 12295
rect 20 12223 18380 12224
rect 20 12219 10251 12223
rect 20 12079 6036 12219
rect 6172 12079 10251 12219
rect 20 12075 10251 12079
rect 10549 12219 18380 12223
rect 10549 12079 12228 12219
rect 12364 12079 18380 12219
rect 10549 12075 18380 12079
rect 20 12074 18380 12075
rect 20 12003 18380 12004
rect 20 11999 5971 12003
rect 20 11859 4488 11999
rect 4624 11859 5971 11999
rect 20 11855 5971 11859
rect 6269 11999 18380 12003
rect 6269 11859 8616 11999
rect 8752 11859 9648 11999
rect 9784 11859 13776 11999
rect 13912 11859 18380 11999
rect 6269 11855 18380 11859
rect 20 11854 18380 11855
rect 20 11783 18380 11784
rect 20 11779 661 11783
rect 899 11779 4341 11783
rect 4579 11779 8021 11783
rect 20 11419 618 11779
rect 899 11419 1134 11779
rect 1270 11419 1650 11779
rect 1786 11419 2166 11779
rect 2302 11419 2682 11779
rect 2818 11419 3198 11779
rect 3334 11419 3714 11779
rect 3850 11419 4230 11779
rect 4579 11419 4746 11779
rect 4882 11419 5262 11779
rect 5398 11419 5778 11779
rect 5914 11419 6294 11779
rect 6430 11419 6810 11779
rect 6946 11419 7326 11779
rect 7462 11419 7842 11779
rect 7978 11419 8021 11779
rect 20 11415 661 11419
rect 899 11415 4341 11419
rect 4579 11415 8021 11419
rect 8259 11779 11701 11783
rect 8259 11419 8358 11779
rect 8494 11419 8874 11779
rect 9010 11419 9390 11779
rect 9526 11419 9906 11779
rect 10042 11419 10422 11779
rect 10558 11419 10938 11779
rect 11074 11419 11454 11779
rect 11590 11419 11701 11779
rect 8259 11415 11701 11419
rect 11939 11779 15381 11783
rect 15619 11779 18380 11783
rect 11939 11419 11970 11779
rect 12106 11419 12486 11779
rect 12622 11419 13002 11779
rect 13138 11419 13518 11779
rect 13654 11419 14034 11779
rect 14170 11419 14550 11779
rect 14686 11419 15066 11779
rect 15202 11419 15381 11779
rect 15718 11419 16098 11779
rect 16234 11419 16614 11779
rect 16750 11419 17130 11779
rect 17266 11419 17646 11779
rect 17782 11419 18380 11779
rect 11939 11415 15381 11419
rect 15619 11415 18380 11419
rect 20 11414 18380 11415
rect 20 11343 18380 11344
rect 20 11339 9651 11343
rect 20 11199 3972 11339
rect 4108 11199 8100 11339
rect 8236 11199 9651 11339
rect 20 11195 9651 11199
rect 9949 11339 18380 11343
rect 9949 11199 10164 11339
rect 10300 11199 14292 11339
rect 14428 11199 18380 11339
rect 9949 11195 18380 11199
rect 20 11194 18380 11195
rect 20 11123 18380 11124
rect 20 11119 6571 11123
rect 6869 11119 18380 11123
rect 20 10979 6552 11119
rect 6869 10979 11712 11119
rect 11848 10979 18380 11119
rect 20 10975 6571 10979
rect 6869 10975 18380 10979
rect 20 10974 18380 10975
rect 20 10903 18380 10904
rect 20 10899 5371 10903
rect 20 10759 2424 10899
rect 2560 10759 5371 10899
rect 20 10755 5371 10759
rect 5669 10899 18380 10903
rect 5669 10759 15840 10899
rect 15976 10759 18380 10899
rect 5669 10755 18380 10759
rect 20 10754 18380 10755
rect 20 10683 18380 10684
rect 20 10679 13931 10683
rect 20 10539 1392 10679
rect 1528 10539 5520 10679
rect 5656 10539 12744 10679
rect 12880 10539 13931 10679
rect 20 10535 13931 10539
rect 14229 10679 18380 10683
rect 14229 10539 16872 10679
rect 17008 10539 18380 10679
rect 14229 10535 18380 10539
rect 20 10534 18380 10535
rect 20 10463 18380 10464
rect 20 10459 12731 10463
rect 20 10319 876 10459
rect 1012 10319 5004 10459
rect 5140 10319 12731 10459
rect 20 10315 12731 10319
rect 13029 10459 18380 10463
rect 13029 10319 13260 10459
rect 13396 10319 17388 10459
rect 17524 10319 18380 10459
rect 13029 10315 18380 10319
rect 20 10314 18380 10315
rect 4634 5846 4681 5910
rect 4745 5846 4751 5910
rect 8314 5846 8361 5910
rect 8425 5846 8431 5910
rect 11994 5846 12041 5910
rect 12105 5846 12111 5910
rect 4634 1224 4801 1288
rect 4865 1224 4871 1288
rect 8314 1224 8481 1288
rect 8545 1224 8551 1288
rect 11994 1224 12161 1288
rect 12225 1224 12231 1288
<< via3 >>
rect 13331 12515 13629 12663
rect 9051 12295 9349 12443
rect 10251 12075 10549 12223
rect 5971 11855 6269 12003
rect 661 11779 899 11783
rect 4341 11779 4579 11783
rect 661 11419 754 11779
rect 754 11419 899 11779
rect 4341 11419 4366 11779
rect 4366 11419 4579 11779
rect 661 11415 899 11419
rect 4341 11415 4579 11419
rect 8021 11415 8259 11783
rect 11701 11415 11939 11783
rect 15381 11779 15619 11783
rect 15381 11419 15582 11779
rect 15582 11419 15619 11779
rect 15381 11415 15619 11419
rect 9651 11195 9949 11343
rect 6571 11119 6869 11123
rect 6571 10979 6688 11119
rect 6688 10979 6869 11119
rect 6571 10975 6869 10979
rect 5371 10755 5669 10903
rect 13931 10535 14229 10683
rect 12731 10315 13029 10463
rect 5971 6147 6269 6545
rect 9651 6147 9949 6545
rect 13331 6147 13629 6545
rect 4681 5846 4745 5910
rect 8361 5846 8425 5910
rect 12041 5846 12105 5910
rect 6571 1525 6869 1923
rect 10251 1525 10549 1923
rect 13931 1525 14229 1923
rect 4801 1224 4865 1288
rect 8481 1224 8545 1288
rect 12161 1224 12225 1288
<< metal4 >>
rect 20 1136 260 12998
rect 340 1136 580 12998
rect 660 11783 900 12998
rect 660 11415 661 11783
rect 899 11415 900 11783
rect 660 -48 900 11415
rect 3700 10198 3940 12998
rect 4020 10198 4260 12998
rect 4340 11783 4580 12998
rect 4340 11415 4341 11783
rect 4579 11415 4580 11783
rect 4340 10198 4580 11415
rect 5370 12698 6270 12998
rect 5370 10903 5670 12698
rect 5370 10755 5371 10903
rect 5669 10755 5670 10903
rect 5370 7846 5670 10755
rect 5970 12003 6270 12004
rect 5970 11855 5971 12003
rect 6269 11855 6270 12003
rect 4680 5910 4746 5911
rect 4680 5846 4681 5910
rect 4745 5846 4746 5910
rect 3700 5576 3940 5846
rect 4020 5576 4260 5846
rect 4340 5576 4580 5846
rect 4680 5845 4746 5846
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1140 4740 5845
rect 5370 3224 5670 7446
rect 5970 6545 6270 11855
rect 5970 6147 5971 6545
rect 6269 6147 6270 6545
rect 5970 6146 6270 6147
rect 6570 11123 6870 11124
rect 6570 10975 6571 11123
rect 6869 10975 6870 11123
rect 6570 1923 6870 10975
rect 7380 10198 7620 12998
rect 7700 10198 7940 12998
rect 8020 11783 8260 12998
rect 8020 11415 8021 11783
rect 8259 11415 8260 11783
rect 8020 10198 8260 11415
rect 9050 12698 9950 12998
rect 9050 12443 9350 12698
rect 9050 12295 9051 12443
rect 9349 12295 9350 12443
rect 9050 7846 9350 12295
rect 10250 12223 10550 12224
rect 10250 12075 10251 12223
rect 10549 12075 10550 12223
rect 9650 11343 9950 11344
rect 9650 11195 9651 11343
rect 9949 11195 9950 11343
rect 8360 5910 8426 5911
rect 8360 5846 8361 5910
rect 8425 5846 8426 5910
rect 7380 5576 7620 5846
rect 7700 5576 7940 5846
rect 8020 5576 8260 5846
rect 8360 5845 8426 5846
rect 6570 1525 6571 1923
rect 6869 1525 6870 1923
rect 6570 1524 6870 1525
rect 4800 1288 4866 1289
rect 4800 1224 4801 1288
rect 4865 1224 4866 1288
rect 4800 1221 4866 1224
rect 4800 1140 4860 1221
rect 7380 1136 7620 1224
rect 7700 1136 7940 1224
rect 8020 -48 8260 1224
rect 8360 1140 8420 5845
rect 9050 3224 9350 7446
rect 9650 6545 9950 11195
rect 9650 6147 9651 6545
rect 9949 6147 9950 6545
rect 9650 6146 9950 6147
rect 10250 1923 10550 12075
rect 11060 10198 11300 12998
rect 11380 10198 11620 12998
rect 11700 11783 11940 12998
rect 11700 11415 11701 11783
rect 11939 11415 11940 11783
rect 11700 10198 11940 11415
rect 13330 12663 13630 12664
rect 13330 12515 13331 12663
rect 13629 12515 13630 12663
rect 12730 10463 13030 10464
rect 12730 10315 12731 10463
rect 13029 10315 13030 10463
rect 12730 7846 13030 10315
rect 12040 5910 12106 5911
rect 12040 5846 12041 5910
rect 12105 5846 12106 5910
rect 11060 5576 11300 5846
rect 11380 5576 11620 5846
rect 11700 5576 11940 5846
rect 12040 5845 12106 5846
rect 10250 1525 10251 1923
rect 10549 1525 10550 1923
rect 10250 1524 10550 1525
rect 8480 1288 8546 1289
rect 8480 1224 8481 1288
rect 8545 1224 8546 1288
rect 8480 1221 8546 1224
rect 8480 1140 8540 1221
rect 11060 1136 11300 1224
rect 11380 1136 11620 1224
rect 11700 -48 11940 1224
rect 12040 1140 12100 5845
rect 12730 3224 13030 7446
rect 13330 6545 13630 12515
rect 13330 6147 13331 6545
rect 13629 6147 13630 6545
rect 13330 6146 13630 6147
rect 13930 10683 14230 10684
rect 13930 10535 13931 10683
rect 14229 10535 14230 10683
rect 13930 1923 14230 10535
rect 13930 1525 13931 1923
rect 14229 1525 14230 1923
rect 13930 1524 14230 1525
rect 12160 1288 12226 1289
rect 12160 1224 12161 1288
rect 12225 1224 12226 1288
rect 12160 1221 12226 1224
rect 12160 1140 12220 1221
rect 14740 1136 14980 13004
rect 15060 1136 15300 13004
rect 15380 11783 15620 12998
rect 15380 11415 15381 11783
rect 15619 11415 15620 11783
rect 15380 -48 15620 11415
use dev_ctrl_b2  dev_ctrl_b2_0
timestamp 1756064790
transform 1 0 11040 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e2  dev_ctrl_e2_0
timestamp 1756064830
transform 1 0 3680 0 1 0
box -38 -48 6868 1140
use dev_ctrl_m2  dev_ctrl_m2_0
timestamp 1756064830
transform 1 0 7360 0 1 0
box -38 -48 6868 1140
use dev_ctrl_p  dev_ctrl_p_0
timestamp 1756676288
transform 1 0 0 0 1 0
box -38 -48 3718 1136
use dev_ctrl_p  dev_ctrl_p_1
timestamp 1756676288
transform 1 0 14720 0 1 0
box -38 -48 3718 1136
use sky130_fd_pr__pfet_g5v0d10v5_L2ZDNS  sky130_fd_pr__pfet_g5v0d10v5_L2ZDNS_0
timestamp 1755863614
transform 1 0 9200 0 1 11599
box -9001 -1047 9001 1047
use tt_asw_3v3  tt_asw_3v3_0
array 0 2 3680 0 1 -4622
timestamp 1756064685
transform 1 0 3680 0 -1 5576
box 0 0 3680 4352
<< end >>
