magic
tech sky130A
magscale 1 2
timestamp 1756676326
<< via3 >>
rect 2291 26763 2589 27161
rect 1691 24311 1989 24609
rect 2291 23711 2589 24009
rect 2291 22141 2589 22539
rect 1691 19689 1989 19987
rect 2291 19089 2589 19387
rect 2291 17519 2589 17917
rect 1691 15067 1989 15365
rect 2291 14467 2589 14765
rect 2291 12897 2589 13295
rect 1691 10445 1989 10743
rect 2291 9845 2589 10143
rect 2291 8275 2589 8673
rect 1691 5823 1989 6121
rect 2291 5223 2589 5521
rect 2291 3653 2589 4051
rect 1691 1201 1989 1499
rect 2291 601 2589 899
<< metal4 >>
rect 2290 27161 2590 27162
rect 2290 26763 2291 27161
rect 2589 26763 2590 27161
rect 1690 24609 1990 25462
rect 1690 24311 1691 24609
rect 1989 24311 1990 24609
rect 1690 24310 1990 24311
rect 2290 24009 2590 26763
rect 2290 23711 2291 24009
rect 2589 23711 2590 24009
rect 2290 23710 2590 23711
rect 2290 22539 2590 22540
rect 2290 22141 2291 22539
rect 2589 22141 2590 22539
rect 1690 19987 1990 20840
rect 1690 19689 1691 19987
rect 1989 19689 1990 19987
rect 1690 19688 1990 19689
rect 2290 19387 2590 22141
rect 2290 19089 2291 19387
rect 2589 19089 2590 19387
rect 2290 19088 2590 19089
rect 2290 17917 2590 17918
rect 2290 17519 2291 17917
rect 2589 17519 2590 17917
rect 1690 15365 1990 16218
rect 1690 15067 1691 15365
rect 1989 15067 1990 15365
rect 1690 15066 1990 15067
rect 2290 14765 2590 17519
rect 2290 14467 2291 14765
rect 2589 14467 2590 14765
rect 2290 14466 2590 14467
rect 2290 13295 2590 13296
rect 2290 12897 2291 13295
rect 2589 12897 2590 13295
rect 1690 10743 1990 11596
rect 1690 10445 1691 10743
rect 1989 10445 1990 10743
rect 1690 10444 1990 10445
rect 2290 10143 2590 12897
rect 2290 9845 2291 10143
rect 2589 9845 2590 10143
rect 2290 9844 2590 9845
rect 2290 8673 2590 8674
rect 2290 8275 2291 8673
rect 2589 8275 2590 8673
rect 1690 6121 1990 6974
rect 1690 5823 1691 6121
rect 1989 5823 1990 6121
rect 1690 5822 1990 5823
rect 2290 5521 2590 8275
rect 2290 5223 2291 5521
rect 2589 5223 2590 5521
rect 2290 5222 2590 5223
rect 2290 4051 2590 4052
rect 2290 3653 2291 4051
rect 2589 3653 2590 4051
rect 1690 1499 1990 2352
rect 1690 1201 1691 1499
rect 1989 1201 1990 1499
rect 1690 1200 1990 1201
rect 2290 899 2590 3653
rect 2290 601 2291 899
rect 2589 601 2590 899
rect 2290 600 2590 601
use asw_col_base  asw_col_base_0
timestamp 1756676326
transform 1 0 0 0 1 0
box -38 0 3718 30910
<< end >>
