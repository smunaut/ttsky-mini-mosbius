magic
tech sky130A
magscale 1 2
timestamp 1756220169
<< nwell >>
rect -1493 -1047 1493 1047
<< mvpmos >>
rect -1235 -750 -1135 750
rect -1077 -750 -977 750
rect -919 -750 -819 750
rect -761 -750 -661 750
rect -603 -750 -503 750
rect -445 -750 -345 750
rect -287 -750 -187 750
rect -129 -750 -29 750
rect 29 -750 129 750
rect 187 -750 287 750
rect 345 -750 445 750
rect 503 -750 603 750
rect 661 -750 761 750
rect 819 -750 919 750
rect 977 -750 1077 750
rect 1135 -750 1235 750
<< mvpdiff >>
rect -1293 738 -1235 750
rect -1293 -738 -1281 738
rect -1247 -738 -1235 738
rect -1293 -750 -1235 -738
rect -1135 738 -1077 750
rect -1135 -738 -1123 738
rect -1089 -738 -1077 738
rect -1135 -750 -1077 -738
rect -977 738 -919 750
rect -977 -738 -965 738
rect -931 -738 -919 738
rect -977 -750 -919 -738
rect -819 738 -761 750
rect -819 -738 -807 738
rect -773 -738 -761 738
rect -819 -750 -761 -738
rect -661 738 -603 750
rect -661 -738 -649 738
rect -615 -738 -603 738
rect -661 -750 -603 -738
rect -503 738 -445 750
rect -503 -738 -491 738
rect -457 -738 -445 738
rect -503 -750 -445 -738
rect -345 738 -287 750
rect -345 -738 -333 738
rect -299 -738 -287 738
rect -345 -750 -287 -738
rect -187 738 -129 750
rect -187 -738 -175 738
rect -141 -738 -129 738
rect -187 -750 -129 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 129 738 187 750
rect 129 -738 141 738
rect 175 -738 187 738
rect 129 -750 187 -738
rect 287 738 345 750
rect 287 -738 299 738
rect 333 -738 345 738
rect 287 -750 345 -738
rect 445 738 503 750
rect 445 -738 457 738
rect 491 -738 503 738
rect 445 -750 503 -738
rect 603 738 661 750
rect 603 -738 615 738
rect 649 -738 661 738
rect 603 -750 661 -738
rect 761 738 819 750
rect 761 -738 773 738
rect 807 -738 819 738
rect 761 -750 819 -738
rect 919 738 977 750
rect 919 -738 931 738
rect 965 -738 977 738
rect 919 -750 977 -738
rect 1077 738 1135 750
rect 1077 -738 1089 738
rect 1123 -738 1135 738
rect 1077 -750 1135 -738
rect 1235 738 1293 750
rect 1235 -738 1247 738
rect 1281 -738 1293 738
rect 1235 -750 1293 -738
<< mvpdiffc >>
rect -1281 -738 -1247 738
rect -1123 -738 -1089 738
rect -965 -738 -931 738
rect -807 -738 -773 738
rect -649 -738 -615 738
rect -491 -738 -457 738
rect -333 -738 -299 738
rect -175 -738 -141 738
rect -17 -738 17 738
rect 141 -738 175 738
rect 299 -738 333 738
rect 457 -738 491 738
rect 615 -738 649 738
rect 773 -738 807 738
rect 931 -738 965 738
rect 1089 -738 1123 738
rect 1247 -738 1281 738
<< mvnsubdiff >>
rect -1427 969 1427 981
rect -1427 935 -1319 969
rect 1319 935 1427 969
rect -1427 923 1427 935
rect -1427 873 -1369 923
rect -1427 -873 -1415 873
rect -1381 -873 -1369 873
rect 1369 873 1427 923
rect -1427 -923 -1369 -873
rect 1369 -873 1381 873
rect 1415 -873 1427 873
rect 1369 -923 1427 -873
rect -1427 -935 1427 -923
rect -1427 -969 -1319 -935
rect 1319 -969 1427 -935
rect -1427 -981 1427 -969
<< mvnsubdiffcont >>
rect -1319 935 1319 969
rect -1415 -873 -1381 873
rect 1381 -873 1415 873
rect -1319 -969 1319 -935
<< poly >>
rect -1235 831 -1135 847
rect -1235 797 -1219 831
rect -1151 797 -1135 831
rect -1235 750 -1135 797
rect -1077 831 -977 847
rect -1077 797 -1061 831
rect -993 797 -977 831
rect -1077 750 -977 797
rect -919 831 -819 847
rect -919 797 -903 831
rect -835 797 -819 831
rect -919 750 -819 797
rect -761 831 -661 847
rect -761 797 -745 831
rect -677 797 -661 831
rect -761 750 -661 797
rect -603 831 -503 847
rect -603 797 -587 831
rect -519 797 -503 831
rect -603 750 -503 797
rect -445 831 -345 847
rect -445 797 -429 831
rect -361 797 -345 831
rect -445 750 -345 797
rect -287 831 -187 847
rect -287 797 -271 831
rect -203 797 -187 831
rect -287 750 -187 797
rect -129 831 -29 847
rect -129 797 -113 831
rect -45 797 -29 831
rect -129 750 -29 797
rect 29 831 129 847
rect 29 797 45 831
rect 113 797 129 831
rect 29 750 129 797
rect 187 831 287 847
rect 187 797 203 831
rect 271 797 287 831
rect 187 750 287 797
rect 345 831 445 847
rect 345 797 361 831
rect 429 797 445 831
rect 345 750 445 797
rect 503 831 603 847
rect 503 797 519 831
rect 587 797 603 831
rect 503 750 603 797
rect 661 831 761 847
rect 661 797 677 831
rect 745 797 761 831
rect 661 750 761 797
rect 819 831 919 847
rect 819 797 835 831
rect 903 797 919 831
rect 819 750 919 797
rect 977 831 1077 847
rect 977 797 993 831
rect 1061 797 1077 831
rect 977 750 1077 797
rect 1135 831 1235 847
rect 1135 797 1151 831
rect 1219 797 1235 831
rect 1135 750 1235 797
rect -1235 -797 -1135 -750
rect -1235 -831 -1219 -797
rect -1151 -831 -1135 -797
rect -1235 -847 -1135 -831
rect -1077 -797 -977 -750
rect -1077 -831 -1061 -797
rect -993 -831 -977 -797
rect -1077 -847 -977 -831
rect -919 -797 -819 -750
rect -919 -831 -903 -797
rect -835 -831 -819 -797
rect -919 -847 -819 -831
rect -761 -797 -661 -750
rect -761 -831 -745 -797
rect -677 -831 -661 -797
rect -761 -847 -661 -831
rect -603 -797 -503 -750
rect -603 -831 -587 -797
rect -519 -831 -503 -797
rect -603 -847 -503 -831
rect -445 -797 -345 -750
rect -445 -831 -429 -797
rect -361 -831 -345 -797
rect -445 -847 -345 -831
rect -287 -797 -187 -750
rect -287 -831 -271 -797
rect -203 -831 -187 -797
rect -287 -847 -187 -831
rect -129 -797 -29 -750
rect -129 -831 -113 -797
rect -45 -831 -29 -797
rect -129 -847 -29 -831
rect 29 -797 129 -750
rect 29 -831 45 -797
rect 113 -831 129 -797
rect 29 -847 129 -831
rect 187 -797 287 -750
rect 187 -831 203 -797
rect 271 -831 287 -797
rect 187 -847 287 -831
rect 345 -797 445 -750
rect 345 -831 361 -797
rect 429 -831 445 -797
rect 345 -847 445 -831
rect 503 -797 603 -750
rect 503 -831 519 -797
rect 587 -831 603 -797
rect 503 -847 603 -831
rect 661 -797 761 -750
rect 661 -831 677 -797
rect 745 -831 761 -797
rect 661 -847 761 -831
rect 819 -797 919 -750
rect 819 -831 835 -797
rect 903 -831 919 -797
rect 819 -847 919 -831
rect 977 -797 1077 -750
rect 977 -831 993 -797
rect 1061 -831 1077 -797
rect 977 -847 1077 -831
rect 1135 -797 1235 -750
rect 1135 -831 1151 -797
rect 1219 -831 1235 -797
rect 1135 -847 1235 -831
<< polycont >>
rect -1219 797 -1151 831
rect -1061 797 -993 831
rect -903 797 -835 831
rect -745 797 -677 831
rect -587 797 -519 831
rect -429 797 -361 831
rect -271 797 -203 831
rect -113 797 -45 831
rect 45 797 113 831
rect 203 797 271 831
rect 361 797 429 831
rect 519 797 587 831
rect 677 797 745 831
rect 835 797 903 831
rect 993 797 1061 831
rect 1151 797 1219 831
rect -1219 -831 -1151 -797
rect -1061 -831 -993 -797
rect -903 -831 -835 -797
rect -745 -831 -677 -797
rect -587 -831 -519 -797
rect -429 -831 -361 -797
rect -271 -831 -203 -797
rect -113 -831 -45 -797
rect 45 -831 113 -797
rect 203 -831 271 -797
rect 361 -831 429 -797
rect 519 -831 587 -797
rect 677 -831 745 -797
rect 835 -831 903 -797
rect 993 -831 1061 -797
rect 1151 -831 1219 -797
<< locali >>
rect -1415 935 -1319 969
rect 1319 935 1415 969
rect -1415 873 -1381 935
rect 1381 873 1415 935
rect -1235 797 -1219 831
rect -1151 797 -1135 831
rect -1077 797 -1061 831
rect -993 797 -977 831
rect -919 797 -903 831
rect -835 797 -819 831
rect -761 797 -745 831
rect -677 797 -661 831
rect -603 797 -587 831
rect -519 797 -503 831
rect -445 797 -429 831
rect -361 797 -345 831
rect -287 797 -271 831
rect -203 797 -187 831
rect -129 797 -113 831
rect -45 797 -29 831
rect 29 797 45 831
rect 113 797 129 831
rect 187 797 203 831
rect 271 797 287 831
rect 345 797 361 831
rect 429 797 445 831
rect 503 797 519 831
rect 587 797 603 831
rect 661 797 677 831
rect 745 797 761 831
rect 819 797 835 831
rect 903 797 919 831
rect 977 797 993 831
rect 1061 797 1077 831
rect 1135 797 1151 831
rect 1219 797 1235 831
rect -1281 738 -1247 754
rect -1281 -754 -1247 -738
rect -1123 738 -1089 754
rect -1123 -754 -1089 -738
rect -965 738 -931 754
rect -965 -754 -931 -738
rect -807 738 -773 754
rect -807 -754 -773 -738
rect -649 738 -615 754
rect -649 -754 -615 -738
rect -491 738 -457 754
rect -491 -754 -457 -738
rect -333 738 -299 754
rect -333 -754 -299 -738
rect -175 738 -141 754
rect -175 -754 -141 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 141 738 175 754
rect 141 -754 175 -738
rect 299 738 333 754
rect 299 -754 333 -738
rect 457 738 491 754
rect 457 -754 491 -738
rect 615 738 649 754
rect 615 -754 649 -738
rect 773 738 807 754
rect 773 -754 807 -738
rect 931 738 965 754
rect 931 -754 965 -738
rect 1089 738 1123 754
rect 1089 -754 1123 -738
rect 1247 738 1281 754
rect 1247 -754 1281 -738
rect -1235 -831 -1219 -797
rect -1151 -831 -1135 -797
rect -1077 -831 -1061 -797
rect -993 -831 -977 -797
rect -919 -831 -903 -797
rect -835 -831 -819 -797
rect -761 -831 -745 -797
rect -677 -831 -661 -797
rect -603 -831 -587 -797
rect -519 -831 -503 -797
rect -445 -831 -429 -797
rect -361 -831 -345 -797
rect -287 -831 -271 -797
rect -203 -831 -187 -797
rect -129 -831 -113 -797
rect -45 -831 -29 -797
rect 29 -831 45 -797
rect 113 -831 129 -797
rect 187 -831 203 -797
rect 271 -831 287 -797
rect 345 -831 361 -797
rect 429 -831 445 -797
rect 503 -831 519 -797
rect 587 -831 603 -797
rect 661 -831 677 -797
rect 745 -831 761 -797
rect 819 -831 835 -797
rect 903 -831 919 -797
rect 977 -831 993 -797
rect 1061 -831 1077 -797
rect 1135 -831 1151 -797
rect 1219 -831 1235 -797
rect -1415 -935 -1381 -873
rect 1381 -935 1415 -873
rect -1415 -969 -1319 -935
rect 1319 -969 1415 -935
<< viali >>
rect -1219 797 -1151 831
rect -1061 797 -993 831
rect -903 797 -835 831
rect -745 797 -677 831
rect -587 797 -519 831
rect -429 797 -361 831
rect -271 797 -203 831
rect -113 797 -45 831
rect 45 797 113 831
rect 203 797 271 831
rect 361 797 429 831
rect 519 797 587 831
rect 677 797 745 831
rect 835 797 903 831
rect 993 797 1061 831
rect 1151 797 1219 831
rect -1281 -738 -1247 738
rect -1123 -738 -1089 738
rect -965 -738 -931 738
rect -807 -738 -773 738
rect -649 -738 -615 738
rect -491 -738 -457 738
rect -333 -738 -299 738
rect -175 -738 -141 738
rect -17 -738 17 738
rect 141 -738 175 738
rect 299 -738 333 738
rect 457 -738 491 738
rect 615 -738 649 738
rect 773 -738 807 738
rect 931 -738 965 738
rect 1089 -738 1123 738
rect 1247 -738 1281 738
rect -1219 -831 -1151 -797
rect -1061 -831 -993 -797
rect -903 -831 -835 -797
rect -745 -831 -677 -797
rect -587 -831 -519 -797
rect -429 -831 -361 -797
rect -271 -831 -203 -797
rect -113 -831 -45 -797
rect 45 -831 113 -797
rect 203 -831 271 -797
rect 361 -831 429 -797
rect 519 -831 587 -797
rect 677 -831 745 -797
rect 835 -831 903 -797
rect 993 -831 1061 -797
rect 1151 -831 1219 -797
<< metal1 >>
rect -1231 831 -1139 837
rect -1231 797 -1219 831
rect -1151 797 -1139 831
rect -1231 791 -1139 797
rect -1073 831 -981 837
rect -1073 797 -1061 831
rect -993 797 -981 831
rect -1073 791 -981 797
rect -915 831 -823 837
rect -915 797 -903 831
rect -835 797 -823 831
rect -915 791 -823 797
rect -757 831 -665 837
rect -757 797 -745 831
rect -677 797 -665 831
rect -757 791 -665 797
rect -599 831 -507 837
rect -599 797 -587 831
rect -519 797 -507 831
rect -599 791 -507 797
rect -441 831 -349 837
rect -441 797 -429 831
rect -361 797 -349 831
rect -441 791 -349 797
rect -283 831 -191 837
rect -283 797 -271 831
rect -203 797 -191 831
rect -283 791 -191 797
rect -125 831 -33 837
rect -125 797 -113 831
rect -45 797 -33 831
rect -125 791 -33 797
rect 33 831 125 837
rect 33 797 45 831
rect 113 797 125 831
rect 33 791 125 797
rect 191 831 283 837
rect 191 797 203 831
rect 271 797 283 831
rect 191 791 283 797
rect 349 831 441 837
rect 349 797 361 831
rect 429 797 441 831
rect 349 791 441 797
rect 507 831 599 837
rect 507 797 519 831
rect 587 797 599 831
rect 507 791 599 797
rect 665 831 757 837
rect 665 797 677 831
rect 745 797 757 831
rect 665 791 757 797
rect 823 831 915 837
rect 823 797 835 831
rect 903 797 915 831
rect 823 791 915 797
rect 981 831 1073 837
rect 981 797 993 831
rect 1061 797 1073 831
rect 981 791 1073 797
rect 1139 831 1231 837
rect 1139 797 1151 831
rect 1219 797 1231 831
rect 1139 791 1231 797
rect -1287 738 -1241 750
rect -1287 -738 -1281 738
rect -1247 -738 -1241 738
rect -1287 -750 -1241 -738
rect -1129 738 -1083 750
rect -1129 -738 -1123 738
rect -1089 -738 -1083 738
rect -1129 -750 -1083 -738
rect -971 738 -925 750
rect -971 -738 -965 738
rect -931 -738 -925 738
rect -971 -750 -925 -738
rect -813 738 -767 750
rect -813 -738 -807 738
rect -773 -738 -767 738
rect -813 -750 -767 -738
rect -655 738 -609 750
rect -655 -738 -649 738
rect -615 -738 -609 738
rect -655 -750 -609 -738
rect -497 738 -451 750
rect -497 -738 -491 738
rect -457 -738 -451 738
rect -497 -750 -451 -738
rect -339 738 -293 750
rect -339 -738 -333 738
rect -299 -738 -293 738
rect -339 -750 -293 -738
rect -181 738 -135 750
rect -181 -738 -175 738
rect -141 -738 -135 738
rect -181 -750 -135 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 135 738 181 750
rect 135 -738 141 738
rect 175 -738 181 738
rect 135 -750 181 -738
rect 293 738 339 750
rect 293 -738 299 738
rect 333 -738 339 738
rect 293 -750 339 -738
rect 451 738 497 750
rect 451 -738 457 738
rect 491 -738 497 738
rect 451 -750 497 -738
rect 609 738 655 750
rect 609 -738 615 738
rect 649 -738 655 738
rect 609 -750 655 -738
rect 767 738 813 750
rect 767 -738 773 738
rect 807 -738 813 738
rect 767 -750 813 -738
rect 925 738 971 750
rect 925 -738 931 738
rect 965 -738 971 738
rect 925 -750 971 -738
rect 1083 738 1129 750
rect 1083 -738 1089 738
rect 1123 -738 1129 738
rect 1083 -750 1129 -738
rect 1241 738 1287 750
rect 1241 -738 1247 738
rect 1281 -738 1287 738
rect 1241 -750 1287 -738
rect -1231 -797 -1139 -791
rect -1231 -831 -1219 -797
rect -1151 -831 -1139 -797
rect -1231 -837 -1139 -831
rect -1073 -797 -981 -791
rect -1073 -831 -1061 -797
rect -993 -831 -981 -797
rect -1073 -837 -981 -831
rect -915 -797 -823 -791
rect -915 -831 -903 -797
rect -835 -831 -823 -797
rect -915 -837 -823 -831
rect -757 -797 -665 -791
rect -757 -831 -745 -797
rect -677 -831 -665 -797
rect -757 -837 -665 -831
rect -599 -797 -507 -791
rect -599 -831 -587 -797
rect -519 -831 -507 -797
rect -599 -837 -507 -831
rect -441 -797 -349 -791
rect -441 -831 -429 -797
rect -361 -831 -349 -797
rect -441 -837 -349 -831
rect -283 -797 -191 -791
rect -283 -831 -271 -797
rect -203 -831 -191 -797
rect -283 -837 -191 -831
rect -125 -797 -33 -791
rect -125 -831 -113 -797
rect -45 -831 -33 -797
rect -125 -837 -33 -831
rect 33 -797 125 -791
rect 33 -831 45 -797
rect 113 -831 125 -797
rect 33 -837 125 -831
rect 191 -797 283 -791
rect 191 -831 203 -797
rect 271 -831 283 -797
rect 191 -837 283 -831
rect 349 -797 441 -791
rect 349 -831 361 -797
rect 429 -831 441 -797
rect 349 -837 441 -831
rect 507 -797 599 -791
rect 507 -831 519 -797
rect 587 -831 599 -797
rect 507 -837 599 -831
rect 665 -797 757 -791
rect 665 -831 677 -797
rect 745 -831 757 -797
rect 665 -837 757 -831
rect 823 -797 915 -791
rect 823 -831 835 -797
rect 903 -831 915 -797
rect 823 -837 915 -831
rect 981 -797 1073 -791
rect 981 -831 993 -797
rect 1061 -831 1073 -797
rect 981 -837 1073 -831
rect 1139 -797 1231 -791
rect 1139 -831 1151 -797
rect 1219 -831 1231 -797
rect 1139 -837 1231 -831
<< labels >>
rlabel mvnsubdiffcont 0 -952 0 -952 0 B
port 1 nsew
rlabel mvpdiffc -1264 0 -1264 0 0 D0
port 2 nsew
rlabel polycont -1185 814 -1185 814 0 G0
port 3 nsew
rlabel mvpdiffc -1106 0 -1106 0 0 S1
port 4 nsew
rlabel polycont -1027 814 -1027 814 0 G1
port 5 nsew
rlabel mvpdiffc -948 0 -948 0 0 D2
port 6 nsew
rlabel polycont -869 814 -869 814 0 G2
port 7 nsew
rlabel mvpdiffc -790 0 -790 0 0 S3
port 8 nsew
rlabel polycont -711 814 -711 814 0 G3
port 9 nsew
rlabel mvpdiffc -632 0 -632 0 0 D4
port 10 nsew
rlabel polycont -553 814 -553 814 0 G4
port 11 nsew
rlabel mvpdiffc -474 0 -474 0 0 S5
port 12 nsew
rlabel polycont -395 814 -395 814 0 G5
port 13 nsew
rlabel mvpdiffc -316 0 -316 0 0 D6
port 14 nsew
rlabel polycont -237 814 -237 814 0 G6
port 15 nsew
rlabel mvpdiffc -158 0 -158 0 0 S7
port 16 nsew
rlabel polycont -79 814 -79 814 0 G7
port 17 nsew
rlabel mvpdiffc 0 0 0 0 0 D8
port 18 nsew
rlabel polycont 79 814 79 814 0 G8
port 19 nsew
rlabel mvpdiffc 158 0 158 0 0 S9
port 20 nsew
rlabel polycont 237 814 237 814 0 G9
port 21 nsew
rlabel mvpdiffc 316 0 316 0 0 D10
port 22 nsew
rlabel polycont 395 814 395 814 0 G10
port 23 nsew
rlabel mvpdiffc 474 0 474 0 0 S11
port 24 nsew
rlabel polycont 553 814 553 814 0 G11
port 25 nsew
rlabel mvpdiffc 632 0 632 0 0 D12
port 26 nsew
rlabel polycont 711 814 711 814 0 G12
port 27 nsew
rlabel mvpdiffc 790 0 790 0 0 S13
port 28 nsew
rlabel polycont 869 814 869 814 0 G13
port 29 nsew
rlabel mvpdiffc 948 0 948 0 0 D14
port 30 nsew
rlabel polycont 1027 814 1027 814 0 G14
port 31 nsew
rlabel mvpdiffc 1106 0 1106 0 0 S15
port 32 nsew
rlabel polycont 1185 814 1185 814 0 G15
port 33 nsew
<< properties >>
string FIXED_BBOX -1398 -952 1398 952
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 0.50 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
