magic
tech sky130A
magscale 1 2
timestamp 1757360412
<< viali >>
rect 215 44507 249 44541
rect 1871 44507 1905 44541
rect 215 43895 249 43929
rect 1871 43895 1905 43929
rect 215 43419 249 43453
rect 1871 43419 1905 43453
rect 97919 41719 97953 41753
rect 98287 41719 98321 41753
rect 8955 1599 8989 1633
rect 9139 1599 9173 1633
rect 9323 1599 9357 1633
rect 7759 1123 7793 1157
rect 9415 1123 9449 1157
<< metal1 >>
rect 200 44498 206 44550
rect 258 44498 264 44550
rect 1856 44498 1862 44550
rect 1914 44498 1920 44550
rect 200 43886 206 43938
rect 258 43886 264 43938
rect 1856 43886 1862 43938
rect 1914 43886 1920 43938
rect 200 43410 206 43462
rect 258 43410 264 43462
rect 1856 43410 1862 43462
rect 1914 43410 1920 43462
rect 2021 42866 2027 42918
rect 2079 42866 2085 42918
rect 1925 41710 1931 41762
rect 1983 41750 1989 41762
rect 97907 41753 97965 41759
rect 97907 41750 97919 41753
rect 1983 41722 2118 41750
rect 97798 41722 97919 41750
rect 1983 41710 1989 41722
rect 97907 41719 97919 41722
rect 97953 41719 97965 41753
rect 97907 41713 97965 41719
rect 98272 41710 98278 41762
rect 98330 41710 98336 41762
rect 8940 1590 8946 1642
rect 8998 1590 9004 1642
rect 9124 1590 9130 1642
rect 9182 1590 9188 1642
rect 9308 1590 9314 1642
rect 9366 1590 9372 1642
rect 7744 1114 7750 1166
rect 7802 1114 7808 1166
rect 9403 1157 9461 1163
rect 9403 1123 9415 1157
rect 9449 1154 9461 1157
rect 9510 1154 9538 1330
rect 9449 1126 9538 1154
rect 9449 1123 9461 1126
rect 9403 1117 9461 1123
<< via1 >>
rect 206 44541 258 44550
rect 206 44507 215 44541
rect 215 44507 249 44541
rect 249 44507 258 44541
rect 206 44498 258 44507
rect 1862 44541 1914 44550
rect 1862 44507 1871 44541
rect 1871 44507 1905 44541
rect 1905 44507 1914 44541
rect 1862 44498 1914 44507
rect 206 43929 258 43938
rect 206 43895 215 43929
rect 215 43895 249 43929
rect 249 43895 258 43929
rect 206 43886 258 43895
rect 1862 43929 1914 43938
rect 1862 43895 1871 43929
rect 1871 43895 1905 43929
rect 1905 43895 1914 43929
rect 1862 43886 1914 43895
rect 206 43453 258 43462
rect 206 43419 215 43453
rect 215 43419 249 43453
rect 249 43419 258 43453
rect 206 43410 258 43419
rect 1862 43453 1914 43462
rect 1862 43419 1871 43453
rect 1871 43419 1905 43453
rect 1905 43419 1914 43453
rect 1862 43410 1914 43419
rect 2027 42909 2079 42918
rect 2027 42875 2036 42909
rect 2036 42875 2070 42909
rect 2070 42875 2079 42909
rect 2027 42866 2079 42875
rect 1931 41710 1983 41762
rect 98278 41753 98330 41762
rect 98278 41719 98287 41753
rect 98287 41719 98321 41753
rect 98321 41719 98330 41753
rect 98278 41710 98330 41719
rect 8946 1633 8998 1642
rect 8946 1599 8955 1633
rect 8955 1599 8989 1633
rect 8989 1599 8998 1633
rect 8946 1590 8998 1599
rect 9130 1633 9182 1642
rect 9130 1599 9139 1633
rect 9139 1599 9173 1633
rect 9173 1599 9182 1633
rect 9130 1590 9182 1599
rect 9314 1633 9366 1642
rect 9314 1599 9323 1633
rect 9323 1599 9357 1633
rect 9357 1599 9366 1633
rect 9314 1590 9366 1599
rect 7750 1157 7802 1166
rect 7750 1123 7759 1157
rect 7759 1123 7793 1157
rect 7793 1123 7802 1157
rect 7750 1114 7802 1123
<< metal2 >>
rect 204 44648 260 44657
rect 204 44550 260 44592
rect 204 44498 206 44550
rect 258 44498 260 44550
rect 204 44492 260 44498
rect 1860 44550 1916 44556
rect 1860 44518 1862 44550
rect 1914 44518 1916 44550
rect 1860 44453 1916 44462
rect 204 44104 260 44113
rect 204 43938 260 44048
rect 204 43886 206 43938
rect 258 43886 260 43938
rect 204 43880 260 43886
rect 1860 43974 1916 43983
rect 1860 43886 1862 43918
rect 1914 43886 1916 43918
rect 1860 43880 1916 43886
rect 204 43560 260 43569
rect 204 43462 260 43504
rect 204 43410 206 43462
rect 258 43410 260 43462
rect 204 43404 260 43410
rect 1860 43462 1916 43468
rect 1860 43430 1862 43462
rect 1914 43430 1916 43462
rect 1860 43365 1916 43374
rect 2025 42920 2081 42929
rect 2025 42855 2081 42864
rect 1929 41764 1985 41773
rect 98383 41762 98392 41764
rect 98272 41710 98278 41762
rect 98330 41710 98392 41762
rect 98383 41708 98392 41710
rect 98448 41708 98457 41764
rect 1929 41699 1985 41708
rect 8944 1644 9000 1653
rect 8944 1579 9000 1588
rect 9128 1644 9184 1653
rect 9128 1579 9184 1588
rect 9312 1644 9368 1653
rect 9312 1579 9368 1588
rect 7748 1168 7804 1177
rect 98383 1166 98392 1168
rect 97594 1114 98392 1166
rect 98383 1112 98392 1114
rect 98448 1112 98457 1168
rect 7748 1103 7804 1112
<< via2 >>
rect 204 44592 260 44648
rect 1860 44498 1862 44518
rect 1862 44498 1914 44518
rect 1914 44498 1916 44518
rect 1860 44462 1916 44498
rect 204 44048 260 44104
rect 1860 43938 1916 43974
rect 1860 43918 1862 43938
rect 1862 43918 1914 43938
rect 1914 43918 1916 43938
rect 204 43504 260 43560
rect 1860 43410 1862 43430
rect 1862 43410 1914 43430
rect 1914 43410 1916 43430
rect 1860 43374 1916 43410
rect 2025 42918 2081 42920
rect 2025 42866 2027 42918
rect 2027 42866 2079 42918
rect 2079 42866 2081 42918
rect 2025 42864 2081 42866
rect 1929 41762 1985 41764
rect 1929 41710 1931 41762
rect 1931 41710 1983 41762
rect 1983 41710 1985 41762
rect 1929 41708 1985 41710
rect 98392 41708 98448 41764
rect 8944 1642 9000 1644
rect 8944 1590 8946 1642
rect 8946 1590 8998 1642
rect 8998 1590 9000 1642
rect 8944 1588 9000 1590
rect 9128 1642 9184 1644
rect 9128 1590 9130 1642
rect 9130 1590 9182 1642
rect 9182 1590 9184 1642
rect 9128 1588 9184 1590
rect 9312 1642 9368 1644
rect 9312 1590 9314 1642
rect 9314 1590 9366 1642
rect 9366 1590 9368 1642
rect 9312 1588 9368 1590
rect 7748 1166 7804 1168
rect 7748 1114 7750 1166
rect 7750 1114 7802 1166
rect 7802 1114 7804 1166
rect 7748 1112 7804 1114
rect 98392 1112 98448 1168
<< metal3 >>
rect 1592 45008 1598 45072
rect 1662 45070 1668 45072
rect 24526 45070 24532 45072
rect 1662 45010 24532 45070
rect 1662 45008 1668 45010
rect 24526 45008 24532 45010
rect 24596 45008 24602 45072
rect 15694 44940 15700 44942
rect 60 44880 15700 44940
rect 60 1170 120 44880
rect 15694 44878 15700 44880
rect 15764 44878 15770 44942
rect 199 44650 265 44653
rect 533 44650 539 44652
rect 199 44648 539 44650
rect 199 44592 204 44648
rect 260 44592 539 44648
rect 199 44590 539 44592
rect 199 44587 265 44590
rect 533 44588 539 44590
rect 603 44588 609 44652
rect 1193 44588 1199 44652
rect 1263 44650 1269 44652
rect 25630 44650 25636 44652
rect 1263 44590 25636 44650
rect 1263 44588 1269 44590
rect 25630 44588 25636 44590
rect 25700 44588 25706 44652
rect 1855 44520 1921 44523
rect 1855 44518 2118 44520
rect 1855 44462 1860 44518
rect 1916 44462 2118 44518
rect 1855 44460 2118 44462
rect 97798 44460 98320 44520
rect 1855 44457 1921 44460
rect 199 44106 265 44109
rect 534 44106 540 44108
rect 199 44104 540 44106
rect 199 44048 204 44104
rect 260 44048 540 44104
rect 199 44046 540 44048
rect 199 44043 265 44046
rect 534 44044 540 44046
rect 604 44044 610 44108
rect 1194 44044 1200 44108
rect 1264 44106 1270 44108
rect 25360 44106 25366 44108
rect 1264 44046 25366 44106
rect 1264 44044 1270 44046
rect 25360 44044 25366 44046
rect 25430 44044 25436 44108
rect 1855 43976 1921 43979
rect 1855 43974 2118 43976
rect 1855 43918 1860 43974
rect 1916 43918 2118 43974
rect 1855 43916 2118 43918
rect 97798 43916 98190 43976
rect 1855 43913 1921 43916
rect 199 43562 265 43565
rect 534 43562 540 43564
rect 199 43560 540 43562
rect 199 43504 204 43560
rect 260 43504 540 43560
rect 199 43502 540 43504
rect 199 43499 265 43502
rect 534 43500 540 43502
rect 604 43500 610 43564
rect 1194 43500 1200 43564
rect 1264 43562 1270 43564
rect 23974 43562 23980 43564
rect 1264 43502 23980 43562
rect 1264 43500 1270 43502
rect 23974 43500 23980 43502
rect 24044 43500 24050 43564
rect 1855 43432 1921 43435
rect 1855 43430 2118 43432
rect 1855 43374 1860 43430
rect 1916 43374 2118 43430
rect 1855 43372 2118 43374
rect 97798 43372 98060 43432
rect 1855 43369 1921 43372
rect 1755 42929 2091 42930
rect 1755 42855 1761 42929
rect 1825 42920 2091 42929
rect 1825 42864 2025 42920
rect 2081 42864 2091 42920
rect 1825 42855 2091 42864
rect 1755 42854 2091 42855
rect 1592 41704 1598 41768
rect 1662 41766 1668 41768
rect 1924 41766 1990 41769
rect 1662 41764 1990 41766
rect 1662 41708 1929 41764
rect 1985 41708 1990 41764
rect 1662 41706 1990 41708
rect 1662 41704 1668 41706
rect 1924 41703 1990 41706
rect 52850 33589 53148 33887
rect 46058 13946 64698 14096
rect 46058 13725 46208 13946
rect 64548 13636 64698 13946
rect 47350 12351 48661 12651
rect 63559 12351 64059 12651
rect 47350 10975 47650 12351
rect 18705 10974 33548 10975
rect 18705 10676 33254 10974
rect 33542 10676 33548 10974
rect 18705 10675 33548 10676
rect 36928 10974 47650 10975
rect 36928 10676 36934 10974
rect 37222 10676 47650 10974
rect 36928 10675 47650 10676
rect 18705 8029 19005 10675
rect 63759 10616 64059 12351
rect 63759 10615 77708 10616
rect 63759 10317 77414 10615
rect 77702 10317 77708 10615
rect 63759 10316 77708 10317
rect 16032 7729 19005 8029
rect 8939 1644 9005 1649
rect 8939 1588 8944 1644
rect 9000 1588 9005 1644
rect 8939 1583 9005 1588
rect 9123 1644 9189 1649
rect 9123 1588 9128 1644
rect 9184 1588 9189 1644
rect 9123 1583 9189 1588
rect 9307 1644 9373 1649
rect 9307 1588 9312 1644
rect 9368 1588 9373 1644
rect 9307 1583 9373 1588
rect 7743 1170 7809 1173
rect 60 1168 7809 1170
rect 60 1112 7748 1168
rect 7804 1112 7809 1168
rect 60 1110 7809 1112
rect 7743 1107 7809 1110
rect 8942 1074 9002 1583
rect 9126 1204 9186 1583
rect 9310 1334 9370 1583
rect 98000 1334 98060 43372
rect 9310 1274 9478 1334
rect 97798 1274 98060 1334
rect 98130 1204 98190 43916
rect 9126 1144 9478 1204
rect 97798 1144 98190 1204
rect 98260 1074 98320 44460
rect 98387 41764 98453 41769
rect 98387 41708 98392 41764
rect 98448 41708 98453 41764
rect 98387 41703 98453 41708
rect 98390 1173 98450 41703
rect 98387 1168 98453 1173
rect 98387 1112 98392 1168
rect 98448 1112 98453 1168
rect 98387 1107 98453 1112
rect 8942 1014 9478 1074
rect 97798 1014 98320 1074
<< via3 >>
rect 1598 45008 1662 45072
rect 24532 45008 24596 45072
rect 15700 44878 15764 44942
rect 539 44588 603 44652
rect 1199 44588 1263 44652
rect 25636 44588 25700 44652
rect 540 44044 604 44108
rect 1200 44044 1264 44108
rect 25366 44044 25430 44108
rect 540 43500 604 43564
rect 1200 43500 1264 43564
rect 23980 43500 24044 43564
rect 1761 42855 1825 42929
rect 1598 41704 1662 41768
rect 19729 38211 20027 38509
rect 63889 37611 64187 37909
rect 67569 33589 67867 33887
rect 5009 32989 5307 33287
rect 52850 28967 53148 29265
rect 8689 28367 8987 28665
rect 12369 24345 12667 24642
rect 56530 23745 56826 24043
rect 47970 15101 48268 15399
rect 59009 14501 59307 14799
rect 32869 11176 33047 11274
rect 33254 10676 33542 10974
rect 36934 10676 37222 10974
rect 77414 10317 77702 10615
<< metal4 >>
rect 1597 45072 1663 45073
rect 1597 45008 1598 45072
rect 1662 45008 1663 45072
rect 3006 45012 3066 45152
rect 3558 45012 3618 45152
rect 4110 45012 4170 45152
rect 4662 45012 4722 45152
rect 5214 45012 5274 45152
rect 5766 45012 5826 45152
rect 6318 45012 6378 45152
rect 6870 45012 6930 45152
rect 7422 45012 7482 45152
rect 7974 45012 8034 45152
rect 8526 45012 8586 45152
rect 9078 45012 9138 45152
rect 9630 45012 9690 45152
rect 10182 45012 10242 45152
rect 10734 45012 10794 45152
rect 11286 45012 11346 45152
rect 11838 45012 11898 45152
rect 12390 45012 12450 45152
rect 12942 45012 13002 45152
rect 13494 45012 13554 45152
rect 14046 45012 14106 45152
rect 14598 45012 14658 45152
rect 15150 45012 15210 45152
rect 1597 45007 1663 45008
rect 538 44652 604 44653
rect 538 44588 539 44652
rect 603 44650 604 44652
rect 1198 44652 1264 44653
rect 1198 44650 1199 44652
rect 603 44590 1199 44650
rect 603 44588 604 44590
rect 538 44587 604 44588
rect 1198 44588 1199 44590
rect 1263 44588 1264 44652
rect 1198 44587 1264 44588
rect 539 44108 605 44109
rect 539 44044 540 44108
rect 604 44106 605 44108
rect 1199 44108 1265 44109
rect 1199 44106 1200 44108
rect 604 44046 1200 44106
rect 604 44044 605 44046
rect 539 44043 605 44044
rect 1199 44044 1200 44046
rect 1264 44044 1265 44108
rect 1199 44043 1265 44044
rect 539 43564 605 43565
rect 539 43500 540 43564
rect 604 43562 605 43564
rect 1199 43564 1265 43565
rect 1199 43562 1200 43564
rect 604 43502 1200 43562
rect 604 43500 605 43502
rect 539 43499 605 43500
rect 1199 43500 1200 43502
rect 1264 43500 1265 43564
rect 1199 43499 1265 43500
rect 1600 41769 1660 45007
rect 1760 44952 15210 45012
rect 1760 42930 1820 44952
rect 15702 44943 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 15699 44942 15765 44943
rect 15699 44878 15700 44942
rect 15764 44878 15765 44942
rect 15699 44877 15765 44878
rect 1760 42929 1826 42930
rect 1760 42855 1761 42929
rect 1825 42855 1826 42929
rect 1760 42854 1826 42855
rect 1597 41768 1663 41769
rect 1597 41704 1598 41768
rect 1662 41704 1663 41768
rect 1597 41703 1663 41704
rect 2138 854 2378 44810
rect 2458 854 2698 44810
rect 2778 854 3018 44810
rect 5008 33287 5308 33288
rect 5008 32989 5009 33287
rect 5307 32989 5308 33287
rect 5008 654 5308 32989
rect 5818 854 6058 44810
rect 6138 854 6378 44810
rect 6458 854 6698 44810
rect 8688 28665 8988 28666
rect 8688 28367 8689 28665
rect 8987 28367 8988 28665
rect 8688 654 8988 28367
rect 9498 854 9738 44810
rect 9818 854 10058 44810
rect 10138 854 10378 44810
rect 12368 24642 12668 24643
rect 12368 24345 12369 24642
rect 12667 24345 12668 24642
rect 12368 654 12668 24345
rect 13178 854 13418 44810
rect 13498 854 13738 44810
rect 13818 854 14058 44810
rect 16858 854 17098 44810
rect 17178 854 17418 44810
rect 17498 854 17738 44810
rect 19728 38509 20028 38510
rect 19728 38211 19729 38509
rect 20027 38211 20028 38509
rect 18528 17252 18828 19722
rect 17978 16952 18828 17252
rect 17978 14800 18278 16952
rect 17978 14500 18828 14800
rect 18528 654 18828 14500
rect 19728 1254 20028 38211
rect 19728 954 20236 1254
rect 19936 654 20236 954
rect 20538 854 20778 44810
rect 20858 854 21098 44810
rect 21178 854 21418 44810
rect 23982 43565 24042 45152
rect 24534 45073 24594 45152
rect 24531 45072 24597 45073
rect 24531 45008 24532 45072
rect 24596 45008 24597 45072
rect 24531 45007 24597 45008
rect 24534 44952 24594 45007
rect 25086 44952 25146 45152
rect 25086 44892 25428 44952
rect 23979 43564 24045 43565
rect 23979 43500 23980 43564
rect 24044 43500 24045 43564
rect 23979 43499 24045 43500
rect 24218 854 24458 44810
rect 24538 854 24778 44810
rect 24858 854 25098 44810
rect 25368 44109 25428 44892
rect 25638 44653 25698 45152
rect 26190 44952 26250 45152
rect 25635 44652 25701 44653
rect 25635 44588 25636 44652
rect 25700 44588 25701 44652
rect 25635 44587 25701 44588
rect 25365 44108 25431 44109
rect 25365 44044 25366 44108
rect 25430 44044 25431 44108
rect 25365 44043 25431 44044
rect 27898 854 28138 44810
rect 28218 854 28458 44810
rect 28538 854 28778 44810
rect 31578 854 31818 44810
rect 31898 854 32138 44810
rect 32218 854 32458 44810
rect 32868 11274 33048 11275
rect 32868 11176 32869 11274
rect 33047 11176 33048 11274
rect 5008 354 8094 654
rect 8688 354 11958 654
rect 12368 354 15822 654
rect 18528 354 19686 654
rect 19936 354 23550 654
rect 32868 380 33048 11176
rect 35258 854 35498 44810
rect 35578 854 35818 44810
rect 35898 854 36138 44810
rect 38938 854 39178 44810
rect 39258 854 39498 44810
rect 39578 854 39818 44810
rect 42618 854 42858 44810
rect 42938 854 43178 44810
rect 43258 854 43498 44810
rect 46298 854 46538 44810
rect 46618 854 46858 44810
rect 46938 854 47178 44810
rect 47969 15399 48269 15400
rect 47969 15101 47970 15399
rect 48268 15101 48269 15399
rect 47969 13900 48269 15101
rect 49978 854 50218 44810
rect 50298 854 50538 44810
rect 50618 854 50858 44810
rect 52849 29265 53149 29266
rect 52849 28967 52850 29265
rect 53148 28967 53149 29265
rect 52849 13900 53149 28967
rect 53658 854 53898 44810
rect 53978 854 54218 44810
rect 54298 854 54538 44810
rect 56529 24043 56827 24044
rect 56529 23745 56530 24043
rect 56826 23745 56827 24043
rect 56529 13900 56827 23745
rect 57338 854 57578 44810
rect 57658 854 57898 44810
rect 57978 854 58218 44810
rect 59008 14799 59308 14800
rect 59008 14501 59009 14799
rect 59307 14501 59308 14799
rect 59008 13900 59308 14501
rect 61018 854 61258 44810
rect 61338 854 61578 44810
rect 61658 854 61898 44810
rect 63888 37909 64188 37910
rect 63888 37611 63889 37909
rect 64187 37611 64188 37909
rect 63888 13900 64188 37611
rect 64698 854 64938 44810
rect 65018 854 65258 44810
rect 65338 854 65578 44810
rect 67568 33887 67868 33888
rect 67568 33589 67569 33887
rect 67867 33589 67868 33887
rect 67568 13900 67868 33589
rect 68378 854 68618 44810
rect 68698 854 68938 44810
rect 69018 854 69258 44810
rect 72058 854 72298 44810
rect 72378 854 72618 44810
rect 72698 854 72938 44810
rect 75738 854 75978 44810
rect 76058 854 76298 44810
rect 76378 854 76618 44810
rect 79418 854 79658 44810
rect 79738 854 79978 44810
rect 80058 854 80298 44810
rect 83098 854 83338 44810
rect 83418 854 83658 44810
rect 83738 854 83978 44810
rect 86778 854 87018 44810
rect 87098 854 87338 44810
rect 87418 854 87658 44810
rect 90458 854 90698 44810
rect 90778 854 91018 44810
rect 91098 854 91338 44810
rect 94138 854 94378 44810
rect 94458 854 94698 44810
rect 94778 854 95018 44810
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 354
rect 11778 0 11958 354
rect 15642 0 15822 354
rect 19506 0 19686 354
rect 23370 0 23550 354
rect 27234 200 33048 380
rect 27234 0 27414 200
<< comment >>
rect -200 45152 98824 45352
rect -200 0 0 45152
rect 98624 0 98824 45152
rect -200 -200 98824 0
use asw_matrix  asw_matrix_0
timestamp 1756676326
transform 1 0 2118 0 1 13900
box -38 0 95718 30910
use dev_ctrl_f  dev_ctrl_f_0
timestamp 1756625277
transform 1 0 94118 0 1 902
box -38 -48 3718 1136
use dev_ctrl_p  dev_ctrl_p_0
timestamp 1756676288
transform 1 0 53638 0 1 902
box -38 -48 3718 1136
use dev_ctrl_p  dev_ctrl_p_2
timestamp 1756676288
transform 1 0 16838 0 1 902
box -38 -48 3718 1136
use dev_nmos_cm  dev_nmos_cm_0
timestamp 1756547599
transform 1 0 31558 0 1 902
box -38 -48 14798 12998
use dev_nmos_dp  dev_nmos_dp_0
timestamp 1756579224
transform 1 0 46278 0 1 902
box -38 -48 10550 12998
use dev_nmos_dual  dev_nmos_dual_0
timestamp 1756547599
transform 1 0 20518 0 1 902
box -1390 -48 17310 13398
use dev_nmos_ota  dev_nmos_ota_0
timestamp 1756710991
transform 1 0 9478 0 1 902
box -1390 -48 7438 12998
use dev_pmos_cm  dev_pmos_cm_0
timestamp 1756676326
transform 1 0 64678 0 1 902
box -38 -48 18438 13004
use dev_pmos_dp  dev_pmos_dp_0
timestamp 1756580837
transform 1 0 57318 0 1 902
box -38 -48 10550 12998
use dev_pmos_dual  dev_pmos_dual_0
timestamp 1756547599
transform 1 0 83078 0 1 902
box -5070 -48 13630 13398
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 97798 0 1 41498
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 186 0 -1 44762
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_1
timestamp 1755005639
transform 1 0 186 0 -1 43674
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_2
timestamp 1755005639
transform 1 0 186 0 1 43674
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_3
timestamp 1755005639
transform -1 0 9478 0 1 902
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  sky130_fd_sc_hd__conb_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 1842 0 1 42586
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 9202 0 -1 1990
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_1
timestamp 1755005639
transform 1 0 9018 0 -1 1990
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  sky130_fd_sc_hd__diode_2_2
timestamp 1755005639
transform 1 0 8834 0 -1 1990
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 2026 0 -1 44762
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1755005639
transform 1 0 2026 0 -1 43674
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1755005639
transform 1 0 2026 0 1 43674
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1755005639
transform 1 0 9386 0 -1 1990
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1755005639
transform 1 0 7546 0 1 902
box -38 -48 130 592
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 2458 854 2698 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 6138 854 6378 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 9818 854 10058 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 13498 854 13738 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 17178 854 17418 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 20858 854 21098 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 24538 854 24778 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 28218 854 28458 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 31898 854 32138 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 35578 854 35818 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 39258 854 39498 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 42938 854 43178 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 46618 854 46858 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 50298 854 50538 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 53978 854 54218 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 57658 854 57898 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 61338 854 61578 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 65018 854 65258 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 68698 854 68938 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 72378 854 72618 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 76058 854 76298 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 79738 854 79978 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 83418 854 83658 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 87098 854 87338 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 90778 854 91018 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 94458 854 94698 44810 0 FreeSans 800 0 0 0 VGND
port 51 nsew ground input
flabel metal4 s 2138 854 2378 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 5818 854 6058 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 9498 854 9738 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 13178 854 13418 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 16858 854 17098 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 20538 854 20778 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 24218 854 24458 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 27898 854 28138 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 31578 854 31818 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 35258 854 35498 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 38938 854 39178 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 42618 854 42858 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 46298 854 46538 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 49978 854 50218 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 53658 854 53898 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 57338 854 57578 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 61018 854 61258 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 64698 854 64938 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 68378 854 68618 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 72058 854 72298 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 75738 854 75978 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 79418 854 79658 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 83098 854 83338 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 86778 854 87018 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 90458 854 90698 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 94138 854 94378 44810 0 FreeSans 800 0 0 0 VDPWR
port 52 nsew power input
flabel metal4 s 2778 854 3018 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 6458 854 6698 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 10138 854 10378 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 13818 854 14058 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 17498 854 17738 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 21178 854 21418 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 24858 854 25098 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 28538 854 28778 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 32218 854 32458 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 35898 854 36138 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 39578 854 39818 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 43258 854 43498 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 46938 854 47178 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 50618 854 50858 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 54298 854 54538 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 57978 854 58218 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 61658 854 61898 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 65338 854 65578 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 69018 854 69258 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 72698 854 72938 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 76378 854 76618 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 80058 854 80298 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 83738 854 83978 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 87418 854 87658 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 91098 854 91338 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
flabel metal4 s 94778 854 95018 44810 0 FreeSans 800 0 0 0 VAPWR
port 53 nsew power input
<< properties >>
string FIXED_BBOX 0 0 98624 45152
<< end >>
