magic
tech sky130A
magscale 1 2
timestamp 1756547599
<< viali >>
rect 4067 12275 6973 12309
rect 3967 10989 4001 12209
rect 5503 10989 5537 12209
rect 7039 10989 7073 12209
rect 4067 10889 6973 10923
<< metal1 >>
rect 4818 12315 4824 12318
rect 3961 12309 4824 12315
rect 6216 12315 6222 12318
rect 6216 12309 7079 12315
rect 3961 12275 4067 12309
rect 6973 12275 7079 12309
rect 3961 12269 4824 12275
rect 3961 12209 4007 12269
rect 4818 12266 4824 12269
rect 6216 12269 7079 12275
rect 6216 12266 6222 12269
rect 3961 10989 3967 12209
rect 4001 10989 4007 12209
rect 5494 12209 5546 12266
rect 5494 12206 5503 12209
rect 5537 12206 5546 12209
rect 4153 12146 4159 12198
rect 5345 12146 5351 12198
rect 4153 12131 5351 12146
rect 4094 12093 4146 12099
rect 4094 11099 4146 11105
rect 4252 12093 4304 12099
rect 4252 11099 4304 11105
rect 4410 12093 4462 12099
rect 4410 11099 4462 11105
rect 4568 12093 4620 12099
rect 4568 11099 4620 11105
rect 4726 12093 4778 12099
rect 4726 11099 4778 11105
rect 4884 12093 4936 12099
rect 4884 11099 4936 11105
rect 5042 12093 5094 12099
rect 5042 11099 5094 11105
rect 5200 12093 5252 12099
rect 5200 11099 5252 11105
rect 5358 12093 5410 12099
rect 5358 11099 5410 11105
rect 4153 11052 5351 11067
rect 4153 11021 4732 11052
rect 4726 11000 4732 11021
rect 5345 11000 5351 11052
rect 3961 10929 4007 10989
rect 7033 12209 7079 12269
rect 5689 12146 5695 12198
rect 6881 12146 6887 12198
rect 5689 12131 6887 12146
rect 5630 12093 5682 12099
rect 5630 11099 5682 11105
rect 5788 12093 5840 12099
rect 5788 11099 5840 11105
rect 5946 12093 5998 12099
rect 5946 11099 5998 11105
rect 6104 12093 6156 12099
rect 6104 11099 6156 11105
rect 6262 12093 6314 12099
rect 6262 11099 6314 11105
rect 6420 12093 6472 12099
rect 6420 11099 6472 11105
rect 6578 12093 6630 12099
rect 6578 11099 6630 11105
rect 6736 12093 6788 12099
rect 6736 11099 6788 11105
rect 6894 12093 6946 12099
rect 6894 11099 6946 11105
rect 5689 11052 6887 11067
rect 5689 11000 5695 11052
rect 6308 11021 6887 11052
rect 6308 11000 6314 11021
rect 5494 10989 5503 10992
rect 5537 10989 5546 10992
rect 5494 10932 5546 10989
rect 7033 10989 7039 12209
rect 7073 10989 7079 12209
rect 4818 10929 4824 10932
rect 3961 10923 4824 10929
rect 6216 10929 6222 10932
rect 7033 10929 7079 10989
rect 6216 10923 7079 10929
rect 3961 10889 4067 10923
rect 6973 10889 7079 10923
rect 3961 10883 4824 10889
rect 4818 10880 4824 10883
rect 6216 10883 7079 10889
rect 6216 10880 6222 10883
<< via1 >>
rect 4824 12309 6216 12318
rect 4824 12275 6216 12309
rect 4824 12266 6216 12275
rect 4159 12146 5345 12198
rect 4094 11105 4146 12093
rect 4252 11105 4304 12093
rect 4410 11105 4462 12093
rect 4568 11105 4620 12093
rect 4726 11105 4778 12093
rect 4884 11105 4936 12093
rect 5042 11105 5094 12093
rect 5200 11105 5252 12093
rect 5358 11105 5410 12093
rect 4732 11000 5345 11052
rect 5494 10992 5503 12206
rect 5503 10992 5537 12206
rect 5537 10992 5546 12206
rect 5695 12146 6881 12198
rect 5630 11105 5682 12093
rect 5788 11105 5840 12093
rect 5946 11105 5998 12093
rect 6104 11105 6156 12093
rect 6262 11105 6314 12093
rect 6420 11105 6472 12093
rect 6578 11105 6630 12093
rect 6736 11105 6788 12093
rect 6894 11105 6946 12093
rect 5695 11000 6308 11052
rect 4824 10923 6216 10932
rect 4824 10889 6216 10923
rect 4824 10880 6216 10889
<< metal2 >>
rect 3958 12294 4754 12299
rect 3958 12204 3967 12294
rect 4745 12204 4754 12294
rect 4818 12266 4824 12318
rect 6216 12266 6222 12318
rect 6286 12294 7082 12299
rect 3958 12198 4754 12204
rect 5494 12206 5546 12266
rect 3958 12146 4159 12198
rect 5345 12146 5351 12198
rect 3958 10932 4010 12146
rect 4092 12094 4148 12103
rect 4092 11795 4094 11804
rect 4146 11795 4148 11804
rect 4252 12093 4304 12103
rect 4210 11694 4252 11703
rect 4368 12094 4504 12103
rect 4368 11795 4410 11804
rect 4304 11694 4346 11703
rect 4210 11495 4252 11504
rect 4094 11095 4146 11105
rect 4304 11495 4346 11504
rect 4252 11095 4304 11105
rect 4462 11795 4504 11804
rect 4568 12093 4620 12103
rect 4410 11095 4462 11105
rect 4526 11194 4568 11203
rect 4684 12094 4820 12103
rect 4684 11795 4726 11804
rect 4620 11194 4662 11203
rect 4778 11795 4820 11804
rect 4884 12093 4936 12103
rect 4842 11394 4884 11403
rect 5000 12094 5136 12103
rect 5000 11795 5042 11804
rect 4936 11394 4978 11403
rect 4842 11235 4884 11244
rect 4726 11095 4778 11105
rect 4936 11235 4978 11244
rect 4884 11095 4936 11105
rect 5094 11795 5136 11804
rect 5200 12093 5252 12103
rect 5158 11694 5200 11703
rect 5356 12094 5412 12103
rect 5356 11795 5358 11804
rect 5252 11694 5294 11703
rect 5158 11495 5200 11504
rect 5042 11095 5094 11105
rect 5252 11495 5294 11504
rect 5200 11095 5252 11105
rect 5410 11795 5412 11804
rect 5358 11095 5410 11105
rect 4526 11035 4662 11044
rect 4726 11000 4732 11052
rect 5345 11000 5351 11052
rect 4726 10932 4778 11000
rect 6286 12204 6295 12294
rect 7073 12204 7082 12294
rect 6286 12198 7082 12204
rect 5689 12146 5695 12198
rect 6881 12146 7082 12198
rect 5628 12094 5684 12103
rect 5628 11795 5630 11804
rect 5682 11795 5684 11804
rect 5788 12093 5840 12103
rect 5746 11694 5788 11703
rect 5904 12094 6040 12103
rect 5904 11795 5946 11804
rect 5840 11694 5882 11703
rect 5746 11495 5788 11504
rect 5630 11095 5682 11105
rect 5840 11495 5882 11504
rect 5788 11095 5840 11105
rect 5998 11795 6040 11804
rect 6104 12093 6156 12103
rect 6062 11394 6104 11403
rect 6220 12094 6356 12103
rect 6220 11795 6262 11804
rect 6156 11394 6198 11403
rect 6062 11235 6104 11244
rect 5946 11095 5998 11105
rect 6156 11235 6198 11244
rect 6104 11095 6156 11105
rect 6314 11795 6356 11804
rect 6420 12093 6472 12103
rect 6262 11095 6314 11105
rect 6378 11194 6420 11203
rect 6536 12094 6672 12103
rect 6536 11795 6578 11804
rect 6472 11194 6514 11203
rect 5689 11000 5695 11052
rect 6308 11000 6314 11052
rect 6630 11795 6672 11804
rect 6736 12093 6788 12103
rect 6694 11694 6736 11703
rect 6892 12094 6948 12103
rect 6892 11795 6894 11804
rect 6788 11694 6830 11703
rect 6694 11495 6736 11504
rect 6578 11095 6630 11105
rect 6788 11495 6830 11504
rect 6736 11095 6788 11105
rect 6946 11795 6948 11804
rect 6894 11095 6946 11105
rect 6378 11035 6514 11044
rect 5494 10932 5546 10992
rect 6262 10932 6314 11000
rect 7030 10932 7082 12146
rect 3958 10880 4778 10932
rect 4818 10880 4824 10932
rect 6216 10880 6222 10932
rect 6262 10880 7082 10932
rect 4818 10837 4827 10880
rect 6213 10837 6222 10880
rect 4818 10832 6222 10837
<< via2 >>
rect 3967 12204 4745 12294
rect 4092 12093 4148 12094
rect 4092 11804 4094 12093
rect 4094 11804 4146 12093
rect 4146 11804 4148 12093
rect 4368 12093 4504 12094
rect 4368 11804 4410 12093
rect 4410 11804 4462 12093
rect 4462 11804 4504 12093
rect 4210 11504 4252 11694
rect 4252 11504 4304 11694
rect 4304 11504 4346 11694
rect 4684 12093 4820 12094
rect 4684 11804 4726 12093
rect 4726 11804 4778 12093
rect 4778 11804 4820 12093
rect 4526 11105 4568 11194
rect 4568 11105 4620 11194
rect 4620 11105 4662 11194
rect 4526 11044 4662 11105
rect 5000 12093 5136 12094
rect 5000 11804 5042 12093
rect 5042 11804 5094 12093
rect 5094 11804 5136 12093
rect 4842 11244 4884 11394
rect 4884 11244 4936 11394
rect 4936 11244 4978 11394
rect 5356 12093 5412 12094
rect 5356 11804 5358 12093
rect 5358 11804 5410 12093
rect 5410 11804 5412 12093
rect 5158 11504 5200 11694
rect 5200 11504 5252 11694
rect 5252 11504 5294 11694
rect 6295 12204 7073 12294
rect 5628 12093 5684 12094
rect 5628 11804 5630 12093
rect 5630 11804 5682 12093
rect 5682 11804 5684 12093
rect 5904 12093 6040 12094
rect 5904 11804 5946 12093
rect 5946 11804 5998 12093
rect 5998 11804 6040 12093
rect 5746 11504 5788 11694
rect 5788 11504 5840 11694
rect 5840 11504 5882 11694
rect 6220 12093 6356 12094
rect 6220 11804 6262 12093
rect 6262 11804 6314 12093
rect 6314 11804 6356 12093
rect 6062 11244 6104 11394
rect 6104 11244 6156 11394
rect 6156 11244 6198 11394
rect 6536 12093 6672 12094
rect 6536 11804 6578 12093
rect 6578 11804 6630 12093
rect 6630 11804 6672 12093
rect 6378 11105 6420 11194
rect 6420 11105 6472 11194
rect 6472 11105 6514 11194
rect 6378 11044 6514 11105
rect 6892 12093 6948 12094
rect 6892 11804 6894 12093
rect 6894 11804 6946 12093
rect 6946 11804 6948 12093
rect 6694 11504 6736 11694
rect 6736 11504 6788 11694
rect 6788 11504 6830 11694
rect 4827 10880 6213 10927
rect 4827 10837 6213 10880
<< metal3 >>
rect 4654 13298 17310 13398
rect -1390 13297 3190 13298
rect -1390 12999 -1384 13297
rect -1096 12999 3190 13297
rect -1390 12998 3190 12999
rect 2890 12099 3190 12998
rect 4654 12299 4754 13298
rect 6982 13197 13630 13198
rect 6982 13098 13336 13197
rect 6982 12299 7082 13098
rect 13330 12999 13336 13098
rect 13624 12999 13630 13197
rect 13330 12998 13630 12999
rect 17010 13197 17310 13298
rect 17010 12999 17016 13197
rect 17304 12999 17310 13197
rect 17010 12998 17310 12999
rect 3958 12294 4754 12299
rect 3958 12204 3967 12294
rect 4745 12204 4754 12294
rect 3958 12199 4754 12204
rect 6286 12294 7082 12299
rect 6286 12204 6295 12294
rect 7073 12204 7082 12294
rect 6286 12199 7082 12204
rect 2890 12098 5417 12099
rect 2890 12094 5113 12098
rect 5411 12094 5417 12098
rect 2890 11804 4092 12094
rect 4148 11804 4368 12094
rect 4504 11804 4684 12094
rect 4820 11804 5000 12094
rect 5412 11804 5417 12094
rect 2890 11800 5113 11804
rect 5411 11800 5417 11804
rect 2890 11799 5417 11800
rect 5623 12098 6953 12099
rect 5623 12094 5971 12098
rect 6269 12094 6953 12098
rect 5623 11804 5628 12094
rect 5684 11804 5904 12094
rect 6356 11804 6536 12094
rect 6672 11804 6892 12094
rect 6948 11804 6953 12094
rect 5623 11800 5971 11804
rect 6269 11800 6953 11804
rect 5623 11799 6953 11800
rect 2885 11698 5299 11699
rect 2885 11500 2891 11698
rect 3189 11694 5299 11698
rect 3189 11504 4210 11694
rect 4346 11504 5158 11694
rect 5294 11504 5299 11694
rect 3189 11500 5299 11504
rect 2885 11499 5299 11500
rect 5741 11698 10555 11699
rect 5741 11694 10251 11698
rect 5741 11504 5746 11694
rect 5882 11504 6694 11694
rect 6830 11504 10251 11694
rect 5741 11500 10251 11504
rect 10549 11500 10555 11698
rect 5741 11499 10555 11500
rect 2285 11498 2595 11499
rect 2285 11300 2291 11498
rect 2589 11399 2595 11498
rect 2589 11394 4983 11399
rect 2589 11300 4842 11394
rect 2285 11299 4842 11300
rect 1685 11298 1995 11299
rect 1685 11100 1691 11298
rect 1989 11199 1995 11298
rect 4837 11244 4842 11299
rect 4978 11244 4983 11394
rect 4837 11239 4983 11244
rect 6057 11398 9955 11399
rect 6057 11394 9651 11398
rect 6057 11244 6062 11394
rect 6198 11299 9651 11394
rect 6198 11244 6203 11299
rect 6057 11239 6203 11244
rect 9645 11200 9651 11299
rect 9949 11200 9955 11398
rect 9645 11199 9955 11200
rect 1989 11194 4667 11199
rect 1989 11100 4526 11194
rect 1685 11099 4526 11100
rect 4521 11044 4526 11099
rect 4662 11044 4667 11194
rect 4521 11039 4667 11044
rect 6373 11198 9355 11199
rect 6373 11194 9051 11198
rect 6373 11044 6378 11194
rect 6514 11099 9051 11194
rect 6514 11044 6519 11099
rect 6373 11039 6519 11044
rect 9045 11000 9051 11099
rect 9349 11000 9355 11198
rect 9045 10999 9355 11000
rect 4020 10931 6222 10932
rect 4020 10833 4026 10931
rect 4254 10927 6222 10931
rect 4254 10837 4827 10927
rect 6213 10837 6222 10927
rect 4254 10833 6222 10837
rect 4020 10832 6222 10833
rect 954 5846 1001 5910
rect 1065 5846 1071 5910
rect 4634 5846 4681 5910
rect 4745 5846 4751 5910
rect 8314 5846 8361 5910
rect 8425 5846 8431 5910
rect 954 1224 1121 1288
rect 1185 1224 1191 1288
rect 4634 1224 4801 1288
rect 4865 1224 4871 1288
rect 8314 1224 8481 1288
rect 8545 1224 8551 1288
<< via3 >>
rect -1384 12999 -1096 13297
rect 13336 12999 13624 13197
rect 17016 12999 17304 13197
rect 5113 12094 5411 12098
rect 5113 11804 5136 12094
rect 5136 11804 5356 12094
rect 5356 11804 5411 12094
rect 5113 11800 5411 11804
rect 5971 12094 6269 12098
rect 5971 11804 6040 12094
rect 6040 11804 6220 12094
rect 6220 11804 6269 12094
rect 5971 11800 6269 11804
rect 2891 11500 3189 11698
rect 10251 11500 10549 11698
rect 2291 11300 2589 11498
rect 1691 11100 1989 11298
rect 9651 11200 9949 11398
rect 9051 11000 9349 11198
rect 4026 10833 4254 10931
rect 4021 7851 4259 8249
rect 2291 6147 2589 6545
rect 5971 6147 6269 6545
rect 9651 6147 9949 6545
rect 1001 5846 1065 5910
rect 4681 5846 4745 5910
rect 8361 5846 8425 5910
rect 4021 3229 4259 3627
rect 2891 1525 3189 1923
rect 6571 1525 6869 1923
rect 10251 1525 10549 1923
rect 1121 1224 1185 1288
rect 4801 1224 4865 1288
rect 8481 1224 8545 1288
<< metal4 >>
rect -1390 13297 -1090 13298
rect -1390 12999 -1384 13297
rect -1096 12999 -1090 13297
rect -1390 12998 -1090 12999
rect 13330 13197 13630 13198
rect 13330 12999 13336 13197
rect 13624 12999 13630 13197
rect 13330 12998 13630 12999
rect 17010 13197 17310 13198
rect 17010 12999 17016 13197
rect 17304 12999 17310 13197
rect 17010 12998 17310 12999
rect 20 10198 260 12998
rect 340 10198 580 12998
rect 660 10198 900 12998
rect 1690 12698 2590 12998
rect 1690 11298 1990 12698
rect 2890 11698 3190 11699
rect 2890 11500 2891 11698
rect 3189 11500 3190 11698
rect 1690 11100 1691 11298
rect 1989 11100 1990 11298
rect 1690 7846 1990 11100
rect 2290 11498 2590 11499
rect 2290 11300 2291 11498
rect 2589 11300 2590 11498
rect 1000 5910 1066 5911
rect 1000 5846 1001 5910
rect 1065 5846 1066 5910
rect 20 5576 260 5846
rect 340 5576 580 5846
rect 660 5576 900 5846
rect 1000 5845 1066 5846
rect 20 1136 260 1224
rect 340 1136 580 1224
rect 660 -48 900 1224
rect 1000 1140 1060 5845
rect 1690 3224 1990 7446
rect 2290 6545 2590 11300
rect 2290 6147 2291 6545
rect 2589 6147 2590 6545
rect 2290 6146 2590 6147
rect 2890 1923 3190 11500
rect 3700 10198 3940 12998
rect 4020 10931 4260 12998
rect 4020 10833 4026 10931
rect 4254 10833 4260 10931
rect 4020 10198 4260 10833
rect 4340 10198 4580 12998
rect 5112 12098 5412 12099
rect 5112 11800 5113 12098
rect 5411 11800 5412 12098
rect 5112 9200 5412 11800
rect 5970 12098 6270 12998
rect 5970 11800 5971 12098
rect 6269 11800 6270 12098
rect 5970 9800 6270 11800
rect 7380 10198 7620 12998
rect 7700 10198 7940 12998
rect 8020 10198 8260 12998
rect 9050 12698 9950 12998
rect 9050 11198 9350 12698
rect 10250 11698 10550 11699
rect 10250 11500 10251 11698
rect 10549 11500 10550 11698
rect 9050 11000 9051 11198
rect 9349 11000 9350 11198
rect 5970 9500 6870 9800
rect 5112 8900 6270 9200
rect 5970 6545 6270 8900
rect 5970 6147 5971 6545
rect 6269 6147 6270 6545
rect 5970 6146 6270 6147
rect 4680 5910 4746 5911
rect 4680 5846 4681 5910
rect 4745 5846 4746 5910
rect 3700 5576 3940 5846
rect 4020 5576 4260 5846
rect 4340 5576 4580 5846
rect 4680 5845 4746 5846
rect 2890 1525 2891 1923
rect 3189 1525 3190 1923
rect 2890 1524 3190 1525
rect 1120 1288 1186 1289
rect 1120 1224 1121 1288
rect 1185 1224 1186 1288
rect 1120 1221 1186 1224
rect 1120 1140 1180 1221
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1140 4740 5845
rect 6570 1923 6870 9500
rect 9050 7846 9350 11000
rect 9650 11398 9950 11399
rect 9650 11200 9651 11398
rect 9949 11200 9950 11398
rect 8360 5910 8426 5911
rect 8360 5846 8361 5910
rect 8425 5846 8426 5910
rect 7380 5576 7620 5846
rect 7700 5576 7940 5846
rect 8020 5576 8260 5846
rect 8360 5845 8426 5846
rect 6570 1525 6571 1923
rect 6869 1525 6870 1923
rect 6570 1524 6870 1525
rect 4800 1288 4866 1289
rect 4800 1224 4801 1288
rect 4865 1224 4866 1288
rect 4800 1221 4866 1224
rect 4800 1140 4860 1221
rect 7380 1136 7620 1224
rect 7700 1136 7940 1224
rect 8020 -48 8260 1224
rect 8360 1140 8420 5845
rect 9050 3224 9350 7446
rect 9650 6545 9950 11200
rect 9650 6147 9651 6545
rect 9949 6147 9950 6545
rect 9650 6146 9950 6147
rect 10250 1923 10550 11500
rect 10250 1525 10251 1923
rect 10549 1525 10550 1923
rect 10250 1524 10550 1525
rect 8480 1288 8546 1289
rect 8480 1224 8481 1288
rect 8545 1224 8546 1288
rect 8480 1221 8546 1224
rect 8480 1140 8540 1221
use dev_ctrl_b2  dev_ctrl_b2_0
timestamp 1756064790
transform 1 0 7360 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e2  dev_ctrl_e2_0
timestamp 1756064830
transform 1 0 0 0 1 0
box -38 -48 6868 1140
use dev_ctrl_m2  dev_ctrl_m2_0
timestamp 1756064830
transform 1 0 3680 0 1 0
box -38 -48 6868 1140
use sky130_fd_pr__nfet_g5v0d10v5_EUEZVQ  sky130_fd_pr__nfet_g5v0d10v5_EUEZVQ_0
timestamp 1756220169
transform 1 0 4752 0 1 11599
box -833 -758 833 758
use sky130_fd_pr__nfet_g5v0d10v5_EUEZVQ  sky130_fd_pr__nfet_g5v0d10v5_EUEZVQ_1
timestamp 1756220169
transform 1 0 6288 0 1 11599
box -833 -758 833 758
use tt_asw_3v3  tt_asw_3v3_0
array 0 2 3680 0 1 -4622
timestamp 1756064685
transform 1 0 0 0 -1 5576
box 0 0 3680 4352
<< properties >>
string FIXED_BBOX 0 0 11040 12998
<< end >>
