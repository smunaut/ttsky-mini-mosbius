magic
tech sky130A
magscale 1 2
timestamp 1756579224
<< viali >>
rect 2363 12275 4997 12309
rect 2263 10989 2297 12209
rect 5063 10989 5097 12209
rect 2363 10889 4997 10923
<< metal1 >>
rect 4020 12315 4026 12318
rect 2257 12309 4026 12315
rect 4254 12315 4260 12318
rect 4254 12309 5103 12315
rect 2257 12275 2363 12309
rect 4997 12275 5103 12309
rect 2257 12269 4026 12275
rect 2257 12209 2303 12269
rect 4020 12266 4026 12269
rect 4254 12269 5103 12275
rect 4254 12266 4260 12269
rect 2257 10989 2263 12209
rect 2297 10989 2303 12209
rect 2469 12227 2521 12233
rect 2627 12227 2679 12233
rect 2541 12131 2607 12177
rect 3101 12227 3153 12233
rect 2857 12131 2923 12177
rect 3259 12227 3311 12233
rect 2785 12080 2837 12086
rect 3173 12131 3239 12177
rect 4049 12227 4101 12233
rect 2943 12080 2995 12086
rect 3489 12131 3555 12177
rect 3417 12080 3469 12086
rect 3575 12080 3627 12086
rect 3805 12131 3871 12177
rect 4207 12227 4259 12233
rect 3733 12080 3785 12086
rect 4121 12131 4187 12177
rect 4681 12227 4733 12233
rect 3891 12080 3943 12086
rect 4437 12131 4503 12177
rect 4839 12227 4891 12233
rect 4365 12080 4417 12086
rect 4753 12131 4819 12177
rect 5057 12209 5103 12269
rect 4523 12080 4575 12086
rect 2390 12043 2442 12049
rect 2390 11149 2442 11155
rect 2548 12043 2600 12049
rect 2548 11149 2600 11155
rect 2706 12043 2758 12049
rect 2706 11149 2758 11155
rect 2864 12043 2916 12049
rect 2864 11149 2916 11155
rect 3022 12043 3074 12049
rect 3022 11149 3074 11155
rect 3180 12043 3232 12049
rect 3180 11149 3232 11155
rect 3338 12043 3390 12049
rect 3338 11149 3390 11155
rect 3496 12043 3548 12049
rect 3496 11149 3548 11155
rect 3654 12043 3706 12049
rect 3654 11149 3706 11155
rect 3812 12043 3864 12049
rect 3812 11149 3864 11155
rect 3970 12043 4022 12049
rect 3970 11149 4022 11155
rect 4128 12043 4180 12049
rect 4128 11149 4180 11155
rect 4286 12043 4338 12049
rect 4286 11149 4338 11155
rect 4444 12043 4496 12049
rect 4444 11149 4496 11155
rect 4602 12043 4654 12049
rect 4602 11149 4654 11155
rect 4760 12043 4812 12049
rect 4760 11149 4812 11155
rect 4918 12043 4970 12049
rect 4918 11149 4970 11155
rect 2469 11112 2521 11118
rect 2627 11112 2679 11118
rect 2541 11021 2607 11067
rect 3101 11112 3153 11118
rect 2257 10929 2303 10989
rect 2857 11021 2923 11067
rect 3259 11112 3311 11118
rect 2785 10965 2837 10971
rect 3173 11021 3239 11067
rect 4049 11112 4101 11118
rect 2943 10965 2995 10971
rect 3489 11021 3555 11067
rect 3417 10965 3469 10971
rect 3575 10965 3627 10971
rect 3805 11021 3871 11067
rect 4207 11112 4259 11118
rect 3733 10965 3785 10971
rect 4121 11021 4187 11067
rect 4681 11112 4733 11118
rect 3891 10965 3943 10971
rect 4437 11021 4503 11067
rect 4839 11112 4891 11118
rect 4365 10965 4417 10971
rect 4753 11021 4819 11067
rect 4523 10965 4575 10971
rect 5057 10989 5063 12209
rect 5097 10989 5103 12209
rect 4020 10929 4026 10932
rect 2257 10923 4026 10929
rect 4254 10929 4260 10932
rect 5057 10929 5103 10989
rect 4254 10923 5103 10929
rect 2257 10889 2363 10923
rect 4997 10889 5103 10923
rect 2257 10883 4026 10889
rect 4020 10880 4026 10883
rect 4254 10883 5103 10889
rect 4254 10880 4260 10883
<< via1 >>
rect 4026 12309 4254 12318
rect 4026 12275 4254 12309
rect 4026 12266 4254 12275
rect 2469 12175 2521 12227
rect 2627 12175 2679 12227
rect 2785 12086 2837 12138
rect 3101 12175 3153 12227
rect 2943 12086 2995 12138
rect 3259 12175 3311 12227
rect 3417 12086 3469 12138
rect 3575 12086 3627 12138
rect 3733 12086 3785 12138
rect 4049 12175 4101 12227
rect 3891 12086 3943 12138
rect 4207 12175 4259 12227
rect 4365 12086 4417 12138
rect 4681 12175 4733 12227
rect 4523 12086 4575 12138
rect 4839 12175 4891 12227
rect 2390 11155 2442 12043
rect 2548 11155 2600 12043
rect 2706 11155 2758 12043
rect 2864 11155 2916 12043
rect 3022 11155 3074 12043
rect 3180 11155 3232 12043
rect 3338 11155 3390 12043
rect 3496 11155 3548 12043
rect 3654 11155 3706 12043
rect 3812 11155 3864 12043
rect 3970 11155 4022 12043
rect 4128 11155 4180 12043
rect 4286 11155 4338 12043
rect 4444 11155 4496 12043
rect 4602 11155 4654 12043
rect 4760 11155 4812 12043
rect 4918 11155 4970 12043
rect 2469 11060 2521 11112
rect 2627 11060 2679 11112
rect 2785 10971 2837 11023
rect 3101 11060 3153 11112
rect 2943 10971 2995 11023
rect 3259 11060 3311 11112
rect 3417 10971 3469 11023
rect 3575 10971 3627 11023
rect 3733 10971 3785 11023
rect 4049 11060 4101 11112
rect 3891 10971 3943 11023
rect 4207 11060 4259 11112
rect 4365 10971 4417 11023
rect 4681 11060 4733 11112
rect 4523 10971 4575 11023
rect 4839 11060 4891 11112
rect 4026 10923 4254 10932
rect 4026 10889 4254 10923
rect 4026 10880 4254 10889
<< metal2 >>
rect 2254 12433 2390 12442
rect 4970 12344 5106 12353
rect 4020 12318 4029 12320
rect 4251 12318 4260 12320
rect 4020 12266 4026 12318
rect 4254 12266 4260 12318
rect 4020 12264 4029 12266
rect 4251 12264 4260 12266
rect 2254 12227 2390 12243
rect 2254 12175 2469 12227
rect 2521 12175 2627 12227
rect 2679 12175 3101 12227
rect 3153 12175 3259 12227
rect 3311 12175 4049 12227
rect 4101 12175 4207 12227
rect 4259 12175 4681 12227
rect 4733 12175 4839 12227
rect 4891 12175 4911 12227
rect 2254 11112 2306 12175
rect 4970 12138 5106 12154
rect 2449 12086 2785 12138
rect 2837 12086 2943 12138
rect 2995 12086 3417 12138
rect 3469 12086 3575 12138
rect 3627 12086 3733 12138
rect 3785 12086 3891 12138
rect 3943 12086 4365 12138
rect 4417 12086 4523 12138
rect 4575 12086 5106 12138
rect 2390 12043 2442 12049
rect 2388 11744 2390 11753
rect 2548 12043 2600 12049
rect 2442 11744 2444 11753
rect 2388 11445 2390 11454
rect 2442 11445 2444 11454
rect 2390 11149 2442 11155
rect 2506 11340 2548 11349
rect 2706 12043 2758 12049
rect 2664 11744 2706 11753
rect 2822 12043 2958 12049
rect 2822 12040 2864 12043
rect 2916 12040 2958 12043
rect 2822 11849 2864 11858
rect 2758 11744 2800 11753
rect 2664 11445 2706 11454
rect 2600 11340 2642 11349
rect 2506 11155 2548 11158
rect 2600 11155 2642 11158
rect 2506 11149 2642 11155
rect 2758 11445 2800 11454
rect 2706 11149 2758 11155
rect 2916 11849 2958 11858
rect 3022 12043 3074 12049
rect 2980 11744 3022 11753
rect 3180 12043 3232 12049
rect 3074 11744 3116 11753
rect 2980 11445 3022 11454
rect 2864 11149 2916 11155
rect 3074 11445 3116 11454
rect 3022 11149 3074 11155
rect 3138 11340 3180 11349
rect 3338 12043 3390 12049
rect 3296 11744 3338 11753
rect 3454 12043 3590 12049
rect 3454 12040 3496 12043
rect 3548 12040 3590 12043
rect 3454 11849 3496 11858
rect 3390 11744 3432 11753
rect 3296 11445 3338 11454
rect 3232 11340 3274 11349
rect 3138 11155 3180 11158
rect 3232 11155 3274 11158
rect 3138 11149 3274 11155
rect 3390 11445 3432 11454
rect 3338 11149 3390 11155
rect 3548 11849 3590 11858
rect 3654 12043 3706 12049
rect 3612 11744 3654 11753
rect 3770 12043 3906 12049
rect 3770 12040 3812 12043
rect 3864 12040 3906 12043
rect 3770 11849 3812 11858
rect 3706 11744 3748 11753
rect 3612 11445 3654 11454
rect 3496 11149 3548 11155
rect 3706 11445 3748 11454
rect 3654 11149 3706 11155
rect 3864 11849 3906 11858
rect 3970 12043 4022 12049
rect 3928 11744 3970 11753
rect 4128 12043 4180 12049
rect 4022 11744 4064 11753
rect 3928 11445 3970 11454
rect 3812 11149 3864 11155
rect 4022 11445 4064 11454
rect 3970 11149 4022 11155
rect 4086 11340 4128 11349
rect 4286 12043 4338 12049
rect 4244 11744 4286 11753
rect 4402 12043 4538 12049
rect 4402 12040 4444 12043
rect 4496 12040 4538 12043
rect 4402 11849 4444 11858
rect 4338 11744 4380 11753
rect 4244 11445 4286 11454
rect 4180 11340 4222 11349
rect 4086 11155 4128 11158
rect 4180 11155 4222 11158
rect 4086 11149 4222 11155
rect 4338 11445 4380 11454
rect 4286 11149 4338 11155
rect 4496 11849 4538 11858
rect 4602 12043 4654 12049
rect 4560 11744 4602 11753
rect 4760 12043 4812 12049
rect 4654 11744 4696 11753
rect 4560 11445 4602 11454
rect 4444 11149 4496 11155
rect 4654 11445 4696 11454
rect 4602 11149 4654 11155
rect 4718 11340 4760 11349
rect 4918 12043 4970 12049
rect 4916 11744 4918 11753
rect 4970 11744 4972 11753
rect 4916 11445 4918 11454
rect 4812 11340 4854 11349
rect 4718 11155 4760 11158
rect 4812 11155 4854 11158
rect 4718 11149 4854 11155
rect 4970 11445 4972 11454
rect 4918 11149 4970 11155
rect 2254 11060 2469 11112
rect 2521 11060 2627 11112
rect 2679 11060 3101 11112
rect 3153 11060 3259 11112
rect 3311 11060 4049 11112
rect 4101 11060 4207 11112
rect 4259 11060 4681 11112
rect 4733 11060 4839 11112
rect 4891 11060 4911 11112
rect 5054 11023 5106 12086
rect 2449 10971 2785 11023
rect 2837 10971 2943 11023
rect 2995 10971 3417 11023
rect 3469 10971 3575 11023
rect 3627 10971 3733 11023
rect 3785 10971 3891 11023
rect 3943 10971 4365 11023
rect 4417 10971 4523 11023
rect 4575 10971 5106 11023
rect 4020 10932 4029 10934
rect 4251 10932 4260 10934
rect 4020 10880 4026 10932
rect 4254 10880 4260 10932
rect 4020 10878 4029 10880
rect 4251 10878 4260 10880
<< via2 >>
rect 2254 12243 2390 12433
rect 4029 12318 4251 12320
rect 4029 12266 4251 12318
rect 4029 12264 4251 12266
rect 4970 12154 5106 12344
rect 2388 11454 2390 11744
rect 2390 11454 2442 11744
rect 2442 11454 2444 11744
rect 2822 11858 2864 12040
rect 2864 11858 2916 12040
rect 2916 11858 2958 12040
rect 2664 11454 2706 11744
rect 2706 11454 2758 11744
rect 2758 11454 2800 11744
rect 2506 11158 2548 11340
rect 2548 11158 2600 11340
rect 2600 11158 2642 11340
rect 2980 11454 3022 11744
rect 3022 11454 3074 11744
rect 3074 11454 3116 11744
rect 3454 11858 3496 12040
rect 3496 11858 3548 12040
rect 3548 11858 3590 12040
rect 3296 11454 3338 11744
rect 3338 11454 3390 11744
rect 3390 11454 3432 11744
rect 3138 11158 3180 11340
rect 3180 11158 3232 11340
rect 3232 11158 3274 11340
rect 3770 11858 3812 12040
rect 3812 11858 3864 12040
rect 3864 11858 3906 12040
rect 3612 11454 3654 11744
rect 3654 11454 3706 11744
rect 3706 11454 3748 11744
rect 3928 11454 3970 11744
rect 3970 11454 4022 11744
rect 4022 11454 4064 11744
rect 4402 11858 4444 12040
rect 4444 11858 4496 12040
rect 4496 11858 4538 12040
rect 4244 11454 4286 11744
rect 4286 11454 4338 11744
rect 4338 11454 4380 11744
rect 4086 11158 4128 11340
rect 4128 11158 4180 11340
rect 4180 11158 4222 11340
rect 4560 11454 4602 11744
rect 4602 11454 4654 11744
rect 4654 11454 4696 11744
rect 4916 11454 4918 11744
rect 4918 11454 4970 11744
rect 4970 11454 4972 11744
rect 4718 11158 4760 11340
rect 4760 11158 4812 11340
rect 4812 11158 4854 11340
rect 4029 10932 4251 10934
rect 4029 10880 4251 10932
rect 4029 10878 4251 10880
<< metal3 >>
rect 2249 12843 2590 12844
rect 2249 12699 2296 12843
rect 2584 12699 2590 12843
rect 2249 12698 2590 12699
rect 2890 12843 5111 12844
rect 2890 12699 2896 12843
rect 3184 12699 5111 12843
rect 2890 12698 5111 12699
rect 2249 12433 2395 12698
rect 2249 12243 2254 12433
rect 2390 12243 2395 12433
rect 4965 12344 5111 12698
rect 4020 12324 4260 12325
rect 4020 12260 4026 12324
rect 4254 12260 4260 12324
rect 4020 12259 4260 12260
rect 2249 12238 2395 12243
rect 4965 12154 4970 12344
rect 5106 12154 5111 12344
rect 4965 12149 5111 12154
rect 2817 12048 9950 12049
rect 2817 12040 9656 12048
rect 2817 11858 2822 12040
rect 2958 11858 3454 12040
rect 3590 11858 3770 12040
rect 3906 11858 4402 12040
rect 4538 11858 9656 12040
rect 2817 11850 9656 11858
rect 9944 11850 9950 12048
rect 2817 11849 9950 11850
rect 2383 11748 4977 11749
rect 2383 11744 2891 11748
rect 3189 11744 4977 11748
rect 2383 11454 2388 11744
rect 2444 11454 2664 11744
rect 2800 11454 2891 11744
rect 3189 11454 3296 11744
rect 3432 11454 3612 11744
rect 3748 11454 3928 11744
rect 4064 11454 4244 11744
rect 4380 11454 4560 11744
rect 4696 11454 4916 11744
rect 4972 11454 4977 11744
rect 2383 11450 2891 11454
rect 3189 11450 4977 11454
rect 2383 11449 4977 11450
rect 2501 11348 6270 11349
rect 2501 11340 5976 11348
rect 2501 11158 2506 11340
rect 2642 11158 3138 11340
rect 3274 11158 4086 11340
rect 4222 11158 4718 11340
rect 4854 11158 5976 11340
rect 2501 11150 5976 11158
rect 6264 11150 6270 11348
rect 2501 11149 6270 11150
rect 4020 10938 4260 10939
rect 4020 10874 4026 10938
rect 4254 10874 4260 10938
rect 4020 10873 4260 10874
rect 7292 8249 10550 8250
rect 7292 7851 10256 8249
rect 10544 7851 10550 8249
rect 7292 7850 10550 7851
rect 954 5846 1001 5910
rect 1065 5846 1071 5910
rect 4634 5846 4681 5910
rect 4745 5846 4751 5910
rect 954 1224 1121 1288
rect 1185 1224 1191 1288
rect 4634 1224 4801 1288
rect 4865 1224 4871 1288
<< via3 >>
rect 2296 12699 2584 12843
rect 2896 12699 3184 12843
rect 4026 12320 4254 12324
rect 4026 12264 4029 12320
rect 4029 12264 4251 12320
rect 4251 12264 4254 12320
rect 4026 12260 4254 12264
rect 9656 11850 9944 12048
rect 2891 11744 3189 11748
rect 2891 11454 2980 11744
rect 2980 11454 3116 11744
rect 3116 11454 3189 11744
rect 2891 11450 3189 11454
rect 5976 11150 6264 11348
rect 4026 10934 4254 10938
rect 4026 10878 4029 10934
rect 4029 10878 4251 10934
rect 4251 10878 4254 10934
rect 4026 10874 4254 10878
rect 341 7851 579 8249
rect 4021 7851 4259 8249
rect 10256 7851 10544 8249
rect 2891 6147 3189 6545
rect 1001 5846 1065 5910
rect 4681 5846 4745 5910
rect 341 3229 579 3627
rect 4021 3229 4259 3627
rect 2291 1525 2589 1923
rect 6571 1525 6869 1923
rect 1121 1224 1185 1288
rect 4801 1224 4865 1288
<< metal4 >>
rect 20 10198 260 12998
rect 340 10198 580 12998
rect 660 10198 900 12998
rect 1691 9200 1990 12998
rect 2290 12843 2590 12998
rect 2290 12699 2296 12843
rect 2584 12699 2590 12843
rect 2290 12698 2590 12699
rect 2890 12843 3190 12998
rect 2890 12699 2896 12843
rect 3184 12699 3190 12843
rect 2890 12698 3190 12699
rect 2890 11748 3190 11749
rect 2890 11450 2891 11748
rect 3189 11450 3190 11748
rect 1691 8900 2590 9200
rect 1000 5910 1066 5911
rect 1000 5846 1001 5910
rect 1065 5846 1066 5910
rect 20 5576 260 5846
rect 340 5576 580 5846
rect 660 5576 900 5846
rect 1000 5845 1066 5846
rect 20 1136 260 1224
rect 340 1136 580 1224
rect 660 -48 900 1224
rect 1000 1140 1060 5845
rect 2290 1923 2590 8900
rect 2890 6545 3190 11450
rect 3700 10198 3940 12998
rect 4020 12324 4260 12998
rect 4020 12260 4026 12324
rect 4254 12260 4260 12324
rect 4020 10938 4260 12260
rect 4020 10874 4026 10938
rect 4254 10874 4260 10938
rect 4020 10198 4260 10874
rect 4340 10198 4580 12998
rect 5970 11348 6270 12998
rect 5970 11150 5976 11348
rect 6264 11150 6270 11348
rect 5970 11149 6270 11150
rect 2890 6147 2891 6545
rect 3189 6147 3190 6545
rect 2890 6146 3190 6147
rect 4680 5910 4746 5911
rect 4680 5846 4681 5910
rect 4745 5846 4746 5910
rect 3700 5576 3940 5846
rect 4020 5576 4260 5846
rect 4340 5576 4580 5846
rect 4680 5845 4746 5846
rect 2290 1525 2291 1923
rect 2589 1525 2590 1923
rect 2290 1524 2590 1525
rect 1120 1288 1186 1289
rect 1120 1224 1121 1288
rect 1185 1224 1186 1288
rect 1120 1221 1186 1224
rect 1120 1140 1180 1221
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1140 4740 5845
rect 6570 1923 6870 12998
rect 9650 12048 9950 12998
rect 9650 11850 9656 12048
rect 9944 11850 9950 12048
rect 9650 11849 9950 11850
rect 10250 8249 10550 12998
rect 10250 7851 10256 8249
rect 10544 7851 10550 8249
rect 10250 7850 10550 7851
rect 6570 1525 6571 1923
rect 6869 1525 6870 1923
rect 6570 1524 6870 1525
rect 4800 1288 4866 1289
rect 4800 1224 4801 1288
rect 4865 1224 4866 1288
rect 4800 1221 4866 1224
rect 4800 1140 4860 1221
use dev_ctrl_b2  dev_ctrl_b2_0
timestamp 1756064790
transform 1 0 3680 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e2  dev_ctrl_e2_0
timestamp 1756064830
transform 1 0 0 0 1 0
box -38 -48 6868 1140
use sky130_fd_pr__nfet_g5v0d10v5_WZKDHM  sky130_fd_pr__nfet_g5v0d10v5_WZKDHM_0
timestamp 1756220169
transform 1 0 3680 0 1 11599
box -1465 -758 1465 758
use tt_asw_3v3  tt_asw_3v3_0
array 0 1 3680 0 1 -4622
timestamp 1756064685
transform 1 0 0 0 -1 5576
box 0 0 3680 4352
<< properties >>
string FIXED_BBOX 0 0 7360 12998
<< end >>
