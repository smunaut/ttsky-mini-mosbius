magic
tech sky130A
magscale 1 2
timestamp 1756547599
<< viali >>
rect 2807 12534 8233 12568
rect 2707 10730 2741 12468
rect 5503 10730 5537 12468
rect 8299 10730 8333 12468
rect 2807 10630 8233 10664
<< metal1 >>
rect 2701 12525 2707 12577
rect 8333 12525 8339 12577
rect 2701 12468 2747 12525
rect 2701 10730 2707 12468
rect 2741 10730 2747 12468
rect 5494 12468 5546 12525
rect 2891 12411 2897 12463
rect 5347 12411 5353 12463
rect 2891 12390 5353 12411
rect 5494 12425 5503 12468
rect 5537 12425 5546 12468
rect 8293 12468 8339 12525
rect 2832 12343 2884 12349
rect 2832 10849 2884 10855
rect 2990 12343 3042 12349
rect 2990 10849 3042 10855
rect 3148 12343 3200 12349
rect 3148 10849 3200 10855
rect 3306 12343 3358 12349
rect 3306 10849 3358 10855
rect 3464 12343 3516 12349
rect 3464 10849 3516 10855
rect 3622 12343 3674 12349
rect 3622 10849 3674 10855
rect 3780 12343 3832 12349
rect 3780 10849 3832 10855
rect 3938 12343 3990 12349
rect 3938 10849 3990 10855
rect 4096 12343 4148 12349
rect 4096 10849 4148 10855
rect 4254 12343 4306 12349
rect 4254 10849 4306 10855
rect 4412 12343 4464 12349
rect 4412 10849 4464 10855
rect 4570 12343 4622 12349
rect 4570 10849 4622 10855
rect 4728 12343 4780 12349
rect 4728 10849 4780 10855
rect 4886 12343 4938 12349
rect 4886 10849 4938 10855
rect 5044 12343 5096 12349
rect 5044 10849 5096 10855
rect 5202 12343 5254 12349
rect 5202 10849 5254 10855
rect 5360 12343 5412 12349
rect 5360 10849 5412 10855
rect 2891 10787 5353 10808
rect 2891 10735 2897 10787
rect 5347 10735 5353 10787
rect 5687 12411 5693 12463
rect 8143 12411 8149 12463
rect 5687 12390 8149 12411
rect 5628 12343 5680 12349
rect 5628 10849 5680 10855
rect 5786 12343 5838 12349
rect 5786 10849 5838 10855
rect 5944 12343 5996 12349
rect 5944 10849 5996 10855
rect 6102 12343 6154 12349
rect 6102 10849 6154 10855
rect 6260 12343 6312 12349
rect 6260 10849 6312 10855
rect 6418 12343 6470 12349
rect 6418 10849 6470 10855
rect 6576 12343 6628 12349
rect 6576 10849 6628 10855
rect 6734 12343 6786 12349
rect 6734 10849 6786 10855
rect 6892 12343 6944 12349
rect 6892 10849 6944 10855
rect 7050 12343 7102 12349
rect 7050 10849 7102 10855
rect 7208 12343 7260 12349
rect 7208 10849 7260 10855
rect 7366 12343 7418 12349
rect 7366 10849 7418 10855
rect 7524 12343 7576 12349
rect 7524 10849 7576 10855
rect 7682 12343 7734 12349
rect 7682 10849 7734 10855
rect 7840 12343 7892 12349
rect 7840 10849 7892 10855
rect 7998 12343 8050 12349
rect 7998 10849 8050 10855
rect 8156 12343 8208 12349
rect 8156 10849 8208 10855
rect 2701 10673 2747 10730
rect 5494 10730 5503 10773
rect 5537 10730 5546 10773
rect 5687 10787 8149 10808
rect 5687 10735 5693 10787
rect 8143 10735 8149 10787
rect 5494 10673 5546 10730
rect 8293 10730 8299 12468
rect 8333 10730 8339 12468
rect 8293 10673 8339 10730
rect 2701 10621 2707 10673
rect 8333 10621 8339 10673
<< via1 >>
rect 2707 12568 8333 12577
rect 2707 12534 2807 12568
rect 2807 12534 8233 12568
rect 8233 12534 8333 12568
rect 2707 12525 8333 12534
rect 2897 12411 5347 12463
rect 2832 10855 2884 12343
rect 2990 10855 3042 12343
rect 3148 10855 3200 12343
rect 3306 10855 3358 12343
rect 3464 10855 3516 12343
rect 3622 10855 3674 12343
rect 3780 10855 3832 12343
rect 3938 10855 3990 12343
rect 4096 10855 4148 12343
rect 4254 10855 4306 12343
rect 4412 10855 4464 12343
rect 4570 10855 4622 12343
rect 4728 10855 4780 12343
rect 4886 10855 4938 12343
rect 5044 10855 5096 12343
rect 5202 10855 5254 12343
rect 5360 10855 5412 12343
rect 2897 10735 5347 10787
rect 5494 10773 5503 12425
rect 5503 10773 5537 12425
rect 5537 10773 5546 12425
rect 5693 12411 8143 12463
rect 5628 10855 5680 12343
rect 5786 10855 5838 12343
rect 5944 10855 5996 12343
rect 6102 10855 6154 12343
rect 6260 10855 6312 12343
rect 6418 10855 6470 12343
rect 6576 10855 6628 12343
rect 6734 10855 6786 12343
rect 6892 10855 6944 12343
rect 7050 10855 7102 12343
rect 7208 10855 7260 12343
rect 7366 10855 7418 12343
rect 7524 10855 7576 12343
rect 7682 10855 7734 12343
rect 7840 10855 7892 12343
rect 7998 10855 8050 12343
rect 8156 10855 8208 12343
rect 5693 10735 8143 10787
rect 2707 10664 8333 10673
rect 2707 10630 2807 10664
rect 2807 10630 8233 10664
rect 8233 10630 8333 10664
rect 2707 10621 8333 10630
<< metal2 >>
rect 2701 12525 2707 12577
rect 8333 12525 8339 12577
rect 2614 12454 2897 12463
rect 2750 12411 2897 12454
rect 5347 12411 5353 12463
rect 5494 12425 5546 12525
rect 2614 12255 2750 12264
rect 2698 10787 2750 12255
rect 2832 12343 2884 12349
rect 2830 11334 2832 11343
rect 2990 12343 3042 12349
rect 2950 11634 2990 11643
rect 3148 12343 3200 12349
rect 3042 11634 3086 11643
rect 2950 11435 2990 11444
rect 2884 11334 2886 11343
rect 2830 11035 2832 11044
rect 2884 11035 2886 11044
rect 2832 10849 2884 10855
rect 3042 11435 3086 11444
rect 3108 11334 3148 11343
rect 3306 12343 3358 12349
rect 3266 11894 3306 11903
rect 3464 12343 3516 12349
rect 3358 11894 3402 11903
rect 3266 11735 3306 11744
rect 3200 11334 3244 11343
rect 3108 11035 3148 11044
rect 2990 10849 3042 10855
rect 3200 11035 3244 11044
rect 3148 10849 3200 10855
rect 3358 11735 3402 11744
rect 3424 11334 3464 11343
rect 3622 12343 3674 12349
rect 3582 12154 3622 12163
rect 3780 12343 3832 12349
rect 3674 12154 3718 12163
rect 3582 11995 3622 12004
rect 3516 11334 3560 11343
rect 3424 11035 3464 11044
rect 3306 10849 3358 10855
rect 3516 11035 3560 11044
rect 3464 10849 3516 10855
rect 3674 11995 3718 12004
rect 3740 11334 3780 11343
rect 3938 12343 3990 12349
rect 3898 11634 3938 11643
rect 4096 12343 4148 12349
rect 3990 11634 4034 11643
rect 3898 11435 3938 11444
rect 3832 11334 3876 11343
rect 3740 11035 3780 11044
rect 3622 10849 3674 10855
rect 3832 11035 3876 11044
rect 3780 10849 3832 10855
rect 3990 11435 4034 11444
rect 4056 11334 4096 11343
rect 4254 12343 4306 12349
rect 4214 11634 4254 11643
rect 4412 12343 4464 12349
rect 4306 11634 4350 11643
rect 4214 11435 4254 11444
rect 4148 11334 4192 11343
rect 4056 11035 4096 11044
rect 3938 10849 3990 10855
rect 4148 11035 4192 11044
rect 4096 10849 4148 10855
rect 4306 11435 4350 11444
rect 4372 11334 4412 11343
rect 4570 12343 4622 12349
rect 4530 12154 4570 12163
rect 4728 12343 4780 12349
rect 4622 12154 4666 12163
rect 4530 11995 4570 12004
rect 4464 11334 4508 11343
rect 4372 11035 4412 11044
rect 4254 10849 4306 10855
rect 4464 11035 4508 11044
rect 4412 10849 4464 10855
rect 4622 11995 4666 12004
rect 4688 11334 4728 11343
rect 4886 12343 4938 12349
rect 4846 11894 4886 11903
rect 5044 12343 5096 12349
rect 4938 11894 4982 11903
rect 4846 11735 4886 11744
rect 4780 11334 4824 11343
rect 4688 11035 4728 11044
rect 4570 10849 4622 10855
rect 4780 11035 4824 11044
rect 4728 10849 4780 10855
rect 4938 11735 4982 11744
rect 5004 11334 5044 11343
rect 5202 12343 5254 12349
rect 5162 11634 5202 11643
rect 5360 12343 5412 12349
rect 5254 11634 5298 11643
rect 5162 11435 5202 11444
rect 5096 11334 5140 11343
rect 5004 11035 5044 11044
rect 4886 10849 4938 10855
rect 5096 11035 5140 11044
rect 5044 10849 5096 10855
rect 5254 11435 5298 11444
rect 5358 11334 5360 11343
rect 5412 11334 5414 11343
rect 5358 11035 5360 11044
rect 5202 10849 5254 10855
rect 5412 11035 5414 11044
rect 5360 10849 5412 10855
rect 2698 10735 2897 10787
rect 5347 10735 5353 10787
rect 5687 12411 5693 12463
rect 8143 12454 8426 12463
rect 8143 12411 8290 12454
rect 5628 12343 5680 12349
rect 5626 11334 5628 11343
rect 5786 12343 5838 12349
rect 5746 11634 5786 11643
rect 5944 12343 5996 12349
rect 5838 11634 5882 11643
rect 5746 11435 5786 11444
rect 5680 11334 5682 11343
rect 5626 11035 5628 11044
rect 5680 11035 5682 11044
rect 5628 10849 5680 10855
rect 5838 11435 5882 11444
rect 5904 11334 5944 11343
rect 6102 12343 6154 12349
rect 6062 11894 6102 11903
rect 6260 12343 6312 12349
rect 6154 11894 6198 11903
rect 6062 11735 6102 11744
rect 5996 11334 6040 11343
rect 5904 11035 5944 11044
rect 5786 10849 5838 10855
rect 5996 11035 6040 11044
rect 5944 10849 5996 10855
rect 6154 11735 6198 11744
rect 6220 11334 6260 11343
rect 6418 12343 6470 12349
rect 6378 12154 6418 12163
rect 6576 12343 6628 12349
rect 6470 12154 6514 12163
rect 6378 11995 6418 12004
rect 6312 11334 6356 11343
rect 6220 11035 6260 11044
rect 6102 10849 6154 10855
rect 6312 11035 6356 11044
rect 6260 10849 6312 10855
rect 6470 11995 6514 12004
rect 6536 11334 6576 11343
rect 6734 12343 6786 12349
rect 6694 11634 6734 11643
rect 6892 12343 6944 12349
rect 6786 11634 6830 11643
rect 6694 11435 6734 11444
rect 6628 11334 6672 11343
rect 6536 11035 6576 11044
rect 6418 10849 6470 10855
rect 6628 11035 6672 11044
rect 6576 10849 6628 10855
rect 6786 11435 6830 11444
rect 6852 11334 6892 11343
rect 7050 12343 7102 12349
rect 7010 11634 7050 11643
rect 7208 12343 7260 12349
rect 7102 11634 7146 11643
rect 7010 11435 7050 11444
rect 6944 11334 6988 11343
rect 6852 11035 6892 11044
rect 6734 10849 6786 10855
rect 6944 11035 6988 11044
rect 6892 10849 6944 10855
rect 7102 11435 7146 11444
rect 7168 11334 7208 11343
rect 7366 12343 7418 12349
rect 7326 12154 7366 12163
rect 7524 12343 7576 12349
rect 7418 12154 7462 12163
rect 7326 11995 7366 12004
rect 7260 11334 7304 11343
rect 7168 11035 7208 11044
rect 7050 10849 7102 10855
rect 7260 11035 7304 11044
rect 7208 10849 7260 10855
rect 7418 11995 7462 12004
rect 7484 11334 7524 11343
rect 7682 12343 7734 12349
rect 7642 11894 7682 11903
rect 7840 12343 7892 12349
rect 7734 11894 7778 11903
rect 7642 11735 7682 11744
rect 7576 11334 7620 11343
rect 7484 11035 7524 11044
rect 7366 10849 7418 10855
rect 7576 11035 7620 11044
rect 7524 10849 7576 10855
rect 7734 11735 7778 11744
rect 7800 11334 7840 11343
rect 7998 12343 8050 12349
rect 7958 11634 7998 11643
rect 8156 12343 8208 12349
rect 8050 11634 8094 11643
rect 7958 11435 7998 11444
rect 7892 11334 7936 11343
rect 7800 11035 7840 11044
rect 7682 10849 7734 10855
rect 7892 11035 7936 11044
rect 7840 10849 7892 10855
rect 8050 11435 8094 11444
rect 8154 11334 8156 11343
rect 8290 12255 8426 12264
rect 8208 11334 8210 11343
rect 8154 11035 8156 11044
rect 7998 10849 8050 10855
rect 8208 11035 8210 11044
rect 8156 10849 8208 10855
rect 8290 10787 8342 12255
rect 5494 10673 5546 10773
rect 5687 10735 5693 10787
rect 8143 10735 8342 10787
rect 2701 10621 2707 10673
rect 8333 10621 8339 10673
rect 4340 10578 4349 10621
rect 6691 10578 6700 10621
rect 4340 10573 6700 10578
<< via2 >>
rect 2614 12264 2750 12454
rect 2950 11444 2990 11634
rect 2990 11444 3042 11634
rect 3042 11444 3086 11634
rect 2830 11044 2832 11334
rect 2832 11044 2884 11334
rect 2884 11044 2886 11334
rect 3266 11744 3306 11894
rect 3306 11744 3358 11894
rect 3358 11744 3402 11894
rect 3108 11044 3148 11334
rect 3148 11044 3200 11334
rect 3200 11044 3244 11334
rect 3582 12004 3622 12154
rect 3622 12004 3674 12154
rect 3674 12004 3718 12154
rect 3424 11044 3464 11334
rect 3464 11044 3516 11334
rect 3516 11044 3560 11334
rect 3898 11444 3938 11634
rect 3938 11444 3990 11634
rect 3990 11444 4034 11634
rect 3740 11044 3780 11334
rect 3780 11044 3832 11334
rect 3832 11044 3876 11334
rect 4214 11444 4254 11634
rect 4254 11444 4306 11634
rect 4306 11444 4350 11634
rect 4056 11044 4096 11334
rect 4096 11044 4148 11334
rect 4148 11044 4192 11334
rect 4530 12004 4570 12154
rect 4570 12004 4622 12154
rect 4622 12004 4666 12154
rect 4372 11044 4412 11334
rect 4412 11044 4464 11334
rect 4464 11044 4508 11334
rect 4846 11744 4886 11894
rect 4886 11744 4938 11894
rect 4938 11744 4982 11894
rect 4688 11044 4728 11334
rect 4728 11044 4780 11334
rect 4780 11044 4824 11334
rect 5162 11444 5202 11634
rect 5202 11444 5254 11634
rect 5254 11444 5298 11634
rect 5004 11044 5044 11334
rect 5044 11044 5096 11334
rect 5096 11044 5140 11334
rect 5358 11044 5360 11334
rect 5360 11044 5412 11334
rect 5412 11044 5414 11334
rect 5746 11444 5786 11634
rect 5786 11444 5838 11634
rect 5838 11444 5882 11634
rect 5626 11044 5628 11334
rect 5628 11044 5680 11334
rect 5680 11044 5682 11334
rect 6062 11744 6102 11894
rect 6102 11744 6154 11894
rect 6154 11744 6198 11894
rect 5904 11044 5944 11334
rect 5944 11044 5996 11334
rect 5996 11044 6040 11334
rect 6378 12004 6418 12154
rect 6418 12004 6470 12154
rect 6470 12004 6514 12154
rect 6220 11044 6260 11334
rect 6260 11044 6312 11334
rect 6312 11044 6356 11334
rect 6694 11444 6734 11634
rect 6734 11444 6786 11634
rect 6786 11444 6830 11634
rect 6536 11044 6576 11334
rect 6576 11044 6628 11334
rect 6628 11044 6672 11334
rect 7010 11444 7050 11634
rect 7050 11444 7102 11634
rect 7102 11444 7146 11634
rect 6852 11044 6892 11334
rect 6892 11044 6944 11334
rect 6944 11044 6988 11334
rect 7326 12004 7366 12154
rect 7366 12004 7418 12154
rect 7418 12004 7462 12154
rect 7168 11044 7208 11334
rect 7208 11044 7260 11334
rect 7260 11044 7304 11334
rect 7642 11744 7682 11894
rect 7682 11744 7734 11894
rect 7734 11744 7778 11894
rect 7484 11044 7524 11334
rect 7524 11044 7576 11334
rect 7576 11044 7620 11334
rect 7958 11444 7998 11634
rect 7998 11444 8050 11634
rect 8050 11444 8094 11634
rect 7800 11044 7840 11334
rect 7840 11044 7892 11334
rect 7892 11044 7936 11334
rect 8290 12264 8426 12454
rect 8154 11044 8156 11334
rect 8156 11044 8208 11334
rect 8208 11044 8210 11334
rect 4349 10621 6691 10668
rect 4349 10578 6691 10621
<< metal3 >>
rect -5070 13298 8408 13398
rect -5070 13197 -4770 13298
rect -5070 12999 -5064 13197
rect -4776 12999 -4770 13197
rect -5070 12998 -4770 12999
rect -1390 13197 2732 13198
rect -1390 12999 -1384 13197
rect -1096 13098 2732 13197
rect -1096 12999 -1090 13098
rect -1390 12998 -1090 12999
rect 2632 12459 2732 13098
rect 8308 12459 8408 13298
rect 10850 13297 13630 13298
rect 10850 12999 13336 13297
rect 13624 12999 13630 13297
rect 10850 12998 13630 12999
rect 2609 12454 2755 12459
rect 2609 12264 2614 12454
rect 2750 12264 2755 12454
rect 2609 12259 2755 12264
rect 8285 12454 8431 12459
rect 8285 12264 8290 12454
rect 8426 12264 8431 12454
rect 8285 12259 8431 12264
rect 1685 12158 4671 12159
rect 1685 12000 1691 12158
rect 1989 12154 4671 12158
rect 1989 12004 3582 12154
rect 3718 12004 4530 12154
rect 4666 12004 4671 12154
rect 1989 12000 4671 12004
rect 1685 11999 4671 12000
rect 6373 12158 9355 12159
rect 6373 12154 9051 12158
rect 6373 12004 6378 12154
rect 6514 12004 7326 12154
rect 7462 12004 9051 12154
rect 6373 12000 9051 12004
rect 9349 12000 9355 12158
rect 6373 11999 9355 12000
rect 2285 11898 4987 11899
rect 2285 11740 2291 11898
rect 2589 11894 4987 11898
rect 2589 11744 3266 11894
rect 3402 11744 4846 11894
rect 4982 11744 4987 11894
rect 2589 11740 4987 11744
rect 2285 11739 4987 11740
rect 6057 11898 9955 11899
rect 6057 11894 9651 11898
rect 6057 11744 6062 11894
rect 6198 11744 7642 11894
rect 7778 11744 9651 11894
rect 6057 11740 9651 11744
rect 9949 11740 9955 11898
rect 6057 11739 9955 11740
rect 2885 11638 5303 11639
rect 2885 11440 2891 11638
rect 3189 11634 5303 11638
rect 3189 11444 3898 11634
rect 4034 11444 4214 11634
rect 4350 11444 5162 11634
rect 5298 11444 5303 11634
rect 3189 11440 5303 11444
rect 2885 11439 5303 11440
rect 5741 11638 10555 11639
rect 5741 11634 10251 11638
rect 5741 11444 5746 11634
rect 5882 11444 6694 11634
rect 6830 11444 7010 11634
rect 7146 11444 7958 11634
rect 8094 11444 10251 11634
rect 5741 11440 10251 11444
rect 10549 11440 10555 11638
rect 5741 11439 10555 11440
rect 10850 11339 11150 12998
rect 2825 11338 5419 11339
rect 2825 11334 5115 11338
rect 5413 11334 5419 11338
rect 2825 11044 2830 11334
rect 2886 11044 3108 11334
rect 3244 11044 3424 11334
rect 3560 11044 3740 11334
rect 3876 11044 4056 11334
rect 4192 11044 4372 11334
rect 4508 11044 4688 11334
rect 4824 11044 5004 11334
rect 5414 11044 5419 11334
rect 2825 11040 5115 11044
rect 5413 11040 5419 11044
rect 2825 11039 5419 11040
rect 5621 11338 11150 11339
rect 5621 11334 6571 11338
rect 6869 11334 11150 11338
rect 5621 11044 5626 11334
rect 5682 11044 5904 11334
rect 6040 11044 6220 11334
rect 6356 11044 6536 11334
rect 6988 11044 7168 11334
rect 7304 11044 7484 11334
rect 7620 11044 7800 11334
rect 7936 11044 8154 11334
rect 8210 11044 11150 11334
rect 5621 11040 6571 11044
rect 6869 11040 11150 11044
rect 5621 11039 11150 11040
rect 4340 10672 6700 10673
rect 4340 10574 4346 10672
rect 4574 10668 6700 10672
rect 6691 10578 6700 10668
rect 4574 10574 6700 10578
rect 4340 10573 6700 10574
rect 954 5846 1001 5910
rect 1065 5846 1071 5910
rect 4634 5846 4681 5910
rect 4745 5846 4751 5910
rect 8314 5846 8361 5910
rect 8425 5846 8431 5910
rect 954 1224 1121 1288
rect 1185 1224 1191 1288
rect 4634 1224 4801 1288
rect 4865 1224 4871 1288
rect 8314 1224 8481 1288
rect 8545 1224 8551 1288
<< via3 >>
rect -5064 12999 -4776 13197
rect -1384 12999 -1096 13197
rect 13336 12999 13624 13297
rect 1691 12000 1989 12158
rect 9051 12000 9349 12158
rect 2291 11740 2589 11898
rect 9651 11740 9949 11898
rect 2891 11634 3189 11638
rect 2891 11444 2950 11634
rect 2950 11444 3086 11634
rect 3086 11444 3189 11634
rect 2891 11440 3189 11444
rect 10251 11440 10549 11638
rect 5115 11334 5413 11338
rect 5115 11044 5140 11334
rect 5140 11044 5358 11334
rect 5358 11044 5413 11334
rect 5115 11040 5413 11044
rect 6571 11334 6869 11338
rect 6571 11044 6672 11334
rect 6672 11044 6852 11334
rect 6852 11044 6869 11334
rect 6571 11040 6869 11044
rect 4346 10668 4574 10672
rect 4346 10578 4349 10668
rect 4349 10578 4574 10668
rect 4346 10574 4574 10578
rect 4341 7851 4579 8249
rect 2291 6147 2589 6545
rect 5971 6147 6269 6545
rect 9651 6147 9949 6545
rect 1001 5846 1065 5910
rect 4681 5846 4745 5910
rect 8361 5846 8425 5910
rect 4341 3229 4579 3627
rect 2891 1525 3189 1923
rect 6571 1525 6869 1923
rect 10251 1525 10549 1923
rect 1121 1224 1185 1288
rect 4801 1224 4865 1288
rect 8481 1224 8545 1288
<< metal4 >>
rect 13330 13297 13630 13298
rect -5070 13197 -4770 13198
rect -5070 12999 -5064 13197
rect -4776 12999 -4770 13197
rect -5070 12998 -4770 12999
rect -1390 13197 -1090 13198
rect -1390 12999 -1384 13197
rect -1096 12999 -1090 13197
rect -1390 12998 -1090 12999
rect 13330 12999 13336 13297
rect 13624 12999 13630 13297
rect 13330 12998 13630 12999
rect 20 10198 260 12998
rect 340 10198 580 12998
rect 660 10198 900 12998
rect 1690 12698 2590 12998
rect 1690 12158 1990 12698
rect 1690 12000 1691 12158
rect 1989 12000 1990 12158
rect 1690 7846 1990 12000
rect 2290 11898 2590 11899
rect 2290 11740 2291 11898
rect 2589 11740 2590 11898
rect 1000 5910 1066 5911
rect 1000 5846 1001 5910
rect 1065 5846 1066 5910
rect 20 5576 260 5846
rect 340 5576 580 5846
rect 660 5576 900 5846
rect 1000 5845 1066 5846
rect 20 1136 260 1224
rect 340 1136 580 1224
rect 660 -48 900 1224
rect 1000 1140 1060 5845
rect 1690 3224 1990 7446
rect 2290 6545 2590 11740
rect 2290 6147 2291 6545
rect 2589 6147 2590 6545
rect 2290 6146 2590 6147
rect 2890 11638 3190 12051
rect 2890 11440 2891 11638
rect 3189 11440 3190 11638
rect 2890 1923 3190 11440
rect 3700 10198 3940 12998
rect 4020 10198 4260 12998
rect 4340 10672 4580 12998
rect 5970 11339 6270 12998
rect 5114 11338 6270 11339
rect 5114 11040 5115 11338
rect 5413 11040 6270 11338
rect 5114 11039 6270 11040
rect 4340 10574 4346 10672
rect 4574 10574 4580 10672
rect 4340 10198 4580 10574
rect 5970 6545 6270 11039
rect 5970 6147 5971 6545
rect 6269 6147 6270 6545
rect 5970 6146 6270 6147
rect 6570 11338 6870 11339
rect 6570 11040 6571 11338
rect 6869 11040 6870 11338
rect 4680 5910 4746 5911
rect 4680 5846 4681 5910
rect 4745 5846 4746 5910
rect 3700 5576 3940 5846
rect 4020 5576 4260 5846
rect 4340 5576 4580 5846
rect 4680 5845 4746 5846
rect 2890 1525 2891 1923
rect 3189 1525 3190 1923
rect 2890 1524 3190 1525
rect 1120 1288 1186 1289
rect 1120 1224 1121 1288
rect 1185 1224 1186 1288
rect 1120 1221 1186 1224
rect 1120 1140 1180 1221
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1140 4740 5845
rect 6570 1923 6870 11040
rect 7380 10198 7620 12998
rect 7700 10198 7940 12998
rect 8020 10198 8260 12998
rect 9050 12698 9950 12998
rect 9050 12158 9350 12698
rect 9050 12000 9051 12158
rect 9349 12000 9350 12158
rect 9050 7846 9350 12000
rect 9650 11898 9950 11899
rect 9650 11740 9651 11898
rect 9949 11740 9950 11898
rect 8360 5910 8426 5911
rect 8360 5846 8361 5910
rect 8425 5846 8426 5910
rect 7380 5576 7620 5846
rect 7700 5576 7940 5846
rect 8020 5576 8260 5846
rect 8360 5845 8426 5846
rect 6570 1525 6571 1923
rect 6869 1525 6870 1923
rect 6570 1524 6870 1525
rect 4800 1288 4866 1289
rect 4800 1224 4801 1288
rect 4865 1224 4866 1288
rect 4800 1221 4866 1224
rect 4800 1140 4860 1221
rect 7380 1136 7620 1224
rect 7700 1136 7940 1224
rect 8020 -48 8260 1224
rect 8360 1140 8420 5845
rect 9050 3224 9350 7446
rect 9650 6545 9950 11740
rect 9650 6147 9651 6545
rect 9949 6147 9950 6545
rect 9650 6146 9950 6147
rect 10250 11638 10550 11639
rect 10250 11440 10251 11638
rect 10549 11440 10550 11638
rect 10250 1923 10550 11440
rect 10250 1525 10251 1923
rect 10549 1525 10550 1923
rect 10250 1524 10550 1525
rect 8480 1288 8546 1289
rect 8480 1224 8481 1288
rect 8545 1224 8546 1288
rect 8480 1221 8546 1224
rect 8480 1140 8540 1221
use dev_ctrl_b2  dev_ctrl_b2_0
timestamp 1756064790
transform 1 0 7360 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e2  dev_ctrl_e2_0
timestamp 1756064830
transform 1 0 0 0 1 0
box -38 -48 6868 1140
use dev_ctrl_m2  dev_ctrl_m2_0
timestamp 1756064830
transform 1 0 3680 0 1 0
box -38 -48 6868 1140
use sky130_fd_pr__pfet_g5v0d10v5_GFVDVM  sky130_fd_pr__pfet_g5v0d10v5_GFVDVM_0
timestamp 1756220169
transform 1 0 4122 0 1 11599
box -1493 -1047 1493 1047
use sky130_fd_pr__pfet_g5v0d10v5_GFVDVM  sky130_fd_pr__pfet_g5v0d10v5_GFVDVM_1
timestamp 1756220169
transform 1 0 6918 0 1 11599
box -1493 -1047 1493 1047
use tt_asw_3v3  tt_asw_3v3_0
array 0 2 3680 0 1 -4622
timestamp 1756064685
transform 1 0 0 0 -1 5576
box 0 0 3680 4352
<< properties >>
string FIXED_BBOX 0 0 11040 12998
<< end >>
