magic
tech sky130A
magscale 1 2
timestamp 1756728921
<< nwell >>
rect -2293 -1047 2293 1047
<< mvpmos >>
rect -2035 -750 -1835 750
rect -1777 -750 -1577 750
rect -1519 -750 -1319 750
rect -1261 -750 -1061 750
rect -1003 -750 -803 750
rect -745 -750 -545 750
rect -487 -750 -287 750
rect -229 -750 -29 750
rect 29 -750 229 750
rect 287 -750 487 750
rect 545 -750 745 750
rect 803 -750 1003 750
rect 1061 -750 1261 750
rect 1319 -750 1519 750
rect 1577 -750 1777 750
rect 1835 -750 2035 750
<< mvpdiff >>
rect -2093 738 -2035 750
rect -2093 -738 -2081 738
rect -2047 -738 -2035 738
rect -2093 -750 -2035 -738
rect -1835 738 -1777 750
rect -1835 -738 -1823 738
rect -1789 -738 -1777 738
rect -1835 -750 -1777 -738
rect -1577 738 -1519 750
rect -1577 -738 -1565 738
rect -1531 -738 -1519 738
rect -1577 -750 -1519 -738
rect -1319 738 -1261 750
rect -1319 -738 -1307 738
rect -1273 -738 -1261 738
rect -1319 -750 -1261 -738
rect -1061 738 -1003 750
rect -1061 -738 -1049 738
rect -1015 -738 -1003 738
rect -1061 -750 -1003 -738
rect -803 738 -745 750
rect -803 -738 -791 738
rect -757 -738 -745 738
rect -803 -750 -745 -738
rect -545 738 -487 750
rect -545 -738 -533 738
rect -499 -738 -487 738
rect -545 -750 -487 -738
rect -287 738 -229 750
rect -287 -738 -275 738
rect -241 -738 -229 738
rect -287 -750 -229 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 229 738 287 750
rect 229 -738 241 738
rect 275 -738 287 738
rect 229 -750 287 -738
rect 487 738 545 750
rect 487 -738 499 738
rect 533 -738 545 738
rect 487 -750 545 -738
rect 745 738 803 750
rect 745 -738 757 738
rect 791 -738 803 738
rect 745 -750 803 -738
rect 1003 738 1061 750
rect 1003 -738 1015 738
rect 1049 -738 1061 738
rect 1003 -750 1061 -738
rect 1261 738 1319 750
rect 1261 -738 1273 738
rect 1307 -738 1319 738
rect 1261 -750 1319 -738
rect 1519 738 1577 750
rect 1519 -738 1531 738
rect 1565 -738 1577 738
rect 1519 -750 1577 -738
rect 1777 738 1835 750
rect 1777 -738 1789 738
rect 1823 -738 1835 738
rect 1777 -750 1835 -738
rect 2035 738 2093 750
rect 2035 -738 2047 738
rect 2081 -738 2093 738
rect 2035 -750 2093 -738
<< mvpdiffc >>
rect -2081 -738 -2047 738
rect -1823 -738 -1789 738
rect -1565 -738 -1531 738
rect -1307 -738 -1273 738
rect -1049 -738 -1015 738
rect -791 -738 -757 738
rect -533 -738 -499 738
rect -275 -738 -241 738
rect -17 -738 17 738
rect 241 -738 275 738
rect 499 -738 533 738
rect 757 -738 791 738
rect 1015 -738 1049 738
rect 1273 -738 1307 738
rect 1531 -738 1565 738
rect 1789 -738 1823 738
rect 2047 -738 2081 738
<< mvnsubdiff >>
rect -2227 969 2227 981
rect -2227 935 -2119 969
rect 2119 935 2227 969
rect -2227 923 2227 935
rect -2227 873 -2169 923
rect -2227 -873 -2215 873
rect -2181 -873 -2169 873
rect 2169 873 2227 923
rect -2227 -923 -2169 -873
rect 2169 -873 2181 873
rect 2215 -873 2227 873
rect 2169 -923 2227 -873
rect -2227 -935 2227 -923
rect -2227 -969 -2119 -935
rect 2119 -969 2227 -935
rect -2227 -981 2227 -969
<< mvnsubdiffcont >>
rect -2119 935 2119 969
rect -2215 -873 -2181 873
rect 2181 -873 2215 873
rect -2119 -969 2119 -935
<< poly >>
rect -2035 831 -1835 847
rect -2035 797 -2019 831
rect -1851 797 -1835 831
rect -2035 750 -1835 797
rect -1777 831 -1577 847
rect -1777 797 -1761 831
rect -1593 797 -1577 831
rect -1777 750 -1577 797
rect -1519 831 -1319 847
rect -1519 797 -1503 831
rect -1335 797 -1319 831
rect -1519 750 -1319 797
rect -1261 831 -1061 847
rect -1261 797 -1245 831
rect -1077 797 -1061 831
rect -1261 750 -1061 797
rect -1003 831 -803 847
rect -1003 797 -987 831
rect -819 797 -803 831
rect -1003 750 -803 797
rect -745 831 -545 847
rect -745 797 -729 831
rect -561 797 -545 831
rect -745 750 -545 797
rect -487 831 -287 847
rect -487 797 -471 831
rect -303 797 -287 831
rect -487 750 -287 797
rect -229 831 -29 847
rect -229 797 -213 831
rect -45 797 -29 831
rect -229 750 -29 797
rect 29 831 229 847
rect 29 797 45 831
rect 213 797 229 831
rect 29 750 229 797
rect 287 831 487 847
rect 287 797 303 831
rect 471 797 487 831
rect 287 750 487 797
rect 545 831 745 847
rect 545 797 561 831
rect 729 797 745 831
rect 545 750 745 797
rect 803 831 1003 847
rect 803 797 819 831
rect 987 797 1003 831
rect 803 750 1003 797
rect 1061 831 1261 847
rect 1061 797 1077 831
rect 1245 797 1261 831
rect 1061 750 1261 797
rect 1319 831 1519 847
rect 1319 797 1335 831
rect 1503 797 1519 831
rect 1319 750 1519 797
rect 1577 831 1777 847
rect 1577 797 1593 831
rect 1761 797 1777 831
rect 1577 750 1777 797
rect 1835 831 2035 847
rect 1835 797 1851 831
rect 2019 797 2035 831
rect 1835 750 2035 797
rect -2035 -797 -1835 -750
rect -2035 -831 -2019 -797
rect -1851 -831 -1835 -797
rect -2035 -847 -1835 -831
rect -1777 -797 -1577 -750
rect -1777 -831 -1761 -797
rect -1593 -831 -1577 -797
rect -1777 -847 -1577 -831
rect -1519 -797 -1319 -750
rect -1519 -831 -1503 -797
rect -1335 -831 -1319 -797
rect -1519 -847 -1319 -831
rect -1261 -797 -1061 -750
rect -1261 -831 -1245 -797
rect -1077 -831 -1061 -797
rect -1261 -847 -1061 -831
rect -1003 -797 -803 -750
rect -1003 -831 -987 -797
rect -819 -831 -803 -797
rect -1003 -847 -803 -831
rect -745 -797 -545 -750
rect -745 -831 -729 -797
rect -561 -831 -545 -797
rect -745 -847 -545 -831
rect -487 -797 -287 -750
rect -487 -831 -471 -797
rect -303 -831 -287 -797
rect -487 -847 -287 -831
rect -229 -797 -29 -750
rect -229 -831 -213 -797
rect -45 -831 -29 -797
rect -229 -847 -29 -831
rect 29 -797 229 -750
rect 29 -831 45 -797
rect 213 -831 229 -797
rect 29 -847 229 -831
rect 287 -797 487 -750
rect 287 -831 303 -797
rect 471 -831 487 -797
rect 287 -847 487 -831
rect 545 -797 745 -750
rect 545 -831 561 -797
rect 729 -831 745 -797
rect 545 -847 745 -831
rect 803 -797 1003 -750
rect 803 -831 819 -797
rect 987 -831 1003 -797
rect 803 -847 1003 -831
rect 1061 -797 1261 -750
rect 1061 -831 1077 -797
rect 1245 -831 1261 -797
rect 1061 -847 1261 -831
rect 1319 -797 1519 -750
rect 1319 -831 1335 -797
rect 1503 -831 1519 -797
rect 1319 -847 1519 -831
rect 1577 -797 1777 -750
rect 1577 -831 1593 -797
rect 1761 -831 1777 -797
rect 1577 -847 1777 -831
rect 1835 -797 2035 -750
rect 1835 -831 1851 -797
rect 2019 -831 2035 -797
rect 1835 -847 2035 -831
<< polycont >>
rect -2019 797 -1851 831
rect -1761 797 -1593 831
rect -1503 797 -1335 831
rect -1245 797 -1077 831
rect -987 797 -819 831
rect -729 797 -561 831
rect -471 797 -303 831
rect -213 797 -45 831
rect 45 797 213 831
rect 303 797 471 831
rect 561 797 729 831
rect 819 797 987 831
rect 1077 797 1245 831
rect 1335 797 1503 831
rect 1593 797 1761 831
rect 1851 797 2019 831
rect -2019 -831 -1851 -797
rect -1761 -831 -1593 -797
rect -1503 -831 -1335 -797
rect -1245 -831 -1077 -797
rect -987 -831 -819 -797
rect -729 -831 -561 -797
rect -471 -831 -303 -797
rect -213 -831 -45 -797
rect 45 -831 213 -797
rect 303 -831 471 -797
rect 561 -831 729 -797
rect 819 -831 987 -797
rect 1077 -831 1245 -797
rect 1335 -831 1503 -797
rect 1593 -831 1761 -797
rect 1851 -831 2019 -797
<< locali >>
rect -2215 935 -2119 969
rect 2119 935 2215 969
rect -2215 873 -2181 935
rect 2181 873 2215 935
rect -2035 797 -2019 831
rect -1851 797 -1835 831
rect -1777 797 -1761 831
rect -1593 797 -1577 831
rect -1519 797 -1503 831
rect -1335 797 -1319 831
rect -1261 797 -1245 831
rect -1077 797 -1061 831
rect -1003 797 -987 831
rect -819 797 -803 831
rect -745 797 -729 831
rect -561 797 -545 831
rect -487 797 -471 831
rect -303 797 -287 831
rect -229 797 -213 831
rect -45 797 -29 831
rect 29 797 45 831
rect 213 797 229 831
rect 287 797 303 831
rect 471 797 487 831
rect 545 797 561 831
rect 729 797 745 831
rect 803 797 819 831
rect 987 797 1003 831
rect 1061 797 1077 831
rect 1245 797 1261 831
rect 1319 797 1335 831
rect 1503 797 1519 831
rect 1577 797 1593 831
rect 1761 797 1777 831
rect 1835 797 1851 831
rect 2019 797 2035 831
rect -2081 738 -2047 754
rect -2081 -754 -2047 -738
rect -1823 738 -1789 754
rect -1823 -754 -1789 -738
rect -1565 738 -1531 754
rect -1565 -754 -1531 -738
rect -1307 738 -1273 754
rect -1307 -754 -1273 -738
rect -1049 738 -1015 754
rect -1049 -754 -1015 -738
rect -791 738 -757 754
rect -791 -754 -757 -738
rect -533 738 -499 754
rect -533 -754 -499 -738
rect -275 738 -241 754
rect -275 -754 -241 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 241 738 275 754
rect 241 -754 275 -738
rect 499 738 533 754
rect 499 -754 533 -738
rect 757 738 791 754
rect 757 -754 791 -738
rect 1015 738 1049 754
rect 1015 -754 1049 -738
rect 1273 738 1307 754
rect 1273 -754 1307 -738
rect 1531 738 1565 754
rect 1531 -754 1565 -738
rect 1789 738 1823 754
rect 1789 -754 1823 -738
rect 2047 738 2081 754
rect 2047 -754 2081 -738
rect -2035 -831 -2019 -797
rect -1851 -831 -1835 -797
rect -1777 -831 -1761 -797
rect -1593 -831 -1577 -797
rect -1519 -831 -1503 -797
rect -1335 -831 -1319 -797
rect -1261 -831 -1245 -797
rect -1077 -831 -1061 -797
rect -1003 -831 -987 -797
rect -819 -831 -803 -797
rect -745 -831 -729 -797
rect -561 -831 -545 -797
rect -487 -831 -471 -797
rect -303 -831 -287 -797
rect -229 -831 -213 -797
rect -45 -831 -29 -797
rect 29 -831 45 -797
rect 213 -831 229 -797
rect 287 -831 303 -797
rect 471 -831 487 -797
rect 545 -831 561 -797
rect 729 -831 745 -797
rect 803 -831 819 -797
rect 987 -831 1003 -797
rect 1061 -831 1077 -797
rect 1245 -831 1261 -797
rect 1319 -831 1335 -797
rect 1503 -831 1519 -797
rect 1577 -831 1593 -797
rect 1761 -831 1777 -797
rect 1835 -831 1851 -797
rect 2019 -831 2035 -797
rect -2215 -935 -2181 -873
rect 2181 -935 2215 -873
rect -2215 -969 -2119 -935
rect 2119 -969 2215 -935
<< viali >>
rect -2019 797 -1851 831
rect -1761 797 -1593 831
rect -1503 797 -1335 831
rect -1245 797 -1077 831
rect -987 797 -819 831
rect -729 797 -561 831
rect -471 797 -303 831
rect -213 797 -45 831
rect 45 797 213 831
rect 303 797 471 831
rect 561 797 729 831
rect 819 797 987 831
rect 1077 797 1245 831
rect 1335 797 1503 831
rect 1593 797 1761 831
rect 1851 797 2019 831
rect -2081 -738 -2047 738
rect -1823 -738 -1789 738
rect -1565 -738 -1531 738
rect -1307 -738 -1273 738
rect -1049 -738 -1015 738
rect -791 -738 -757 738
rect -533 -738 -499 738
rect -275 -738 -241 738
rect -17 -738 17 738
rect 241 -738 275 738
rect 499 -738 533 738
rect 757 -738 791 738
rect 1015 -738 1049 738
rect 1273 -738 1307 738
rect 1531 -738 1565 738
rect 1789 -738 1823 738
rect 2047 -738 2081 738
rect -2019 -831 -1851 -797
rect -1761 -831 -1593 -797
rect -1503 -831 -1335 -797
rect -1245 -831 -1077 -797
rect -987 -831 -819 -797
rect -729 -831 -561 -797
rect -471 -831 -303 -797
rect -213 -831 -45 -797
rect 45 -831 213 -797
rect 303 -831 471 -797
rect 561 -831 729 -797
rect 819 -831 987 -797
rect 1077 -831 1245 -797
rect 1335 -831 1503 -797
rect 1593 -831 1761 -797
rect 1851 -831 2019 -797
<< metal1 >>
rect -2031 831 -1839 837
rect -2031 797 -2019 831
rect -1851 797 -1839 831
rect -2031 791 -1839 797
rect -1773 831 -1581 837
rect -1773 797 -1761 831
rect -1593 797 -1581 831
rect -1773 791 -1581 797
rect -1515 831 -1323 837
rect -1515 797 -1503 831
rect -1335 797 -1323 831
rect -1515 791 -1323 797
rect -1257 831 -1065 837
rect -1257 797 -1245 831
rect -1077 797 -1065 831
rect -1257 791 -1065 797
rect -999 831 -807 837
rect -999 797 -987 831
rect -819 797 -807 831
rect -999 791 -807 797
rect -741 831 -549 837
rect -741 797 -729 831
rect -561 797 -549 831
rect -741 791 -549 797
rect -483 831 -291 837
rect -483 797 -471 831
rect -303 797 -291 831
rect -483 791 -291 797
rect -225 831 -33 837
rect -225 797 -213 831
rect -45 797 -33 831
rect -225 791 -33 797
rect 33 831 225 837
rect 33 797 45 831
rect 213 797 225 831
rect 33 791 225 797
rect 291 831 483 837
rect 291 797 303 831
rect 471 797 483 831
rect 291 791 483 797
rect 549 831 741 837
rect 549 797 561 831
rect 729 797 741 831
rect 549 791 741 797
rect 807 831 999 837
rect 807 797 819 831
rect 987 797 999 831
rect 807 791 999 797
rect 1065 831 1257 837
rect 1065 797 1077 831
rect 1245 797 1257 831
rect 1065 791 1257 797
rect 1323 831 1515 837
rect 1323 797 1335 831
rect 1503 797 1515 831
rect 1323 791 1515 797
rect 1581 831 1773 837
rect 1581 797 1593 831
rect 1761 797 1773 831
rect 1581 791 1773 797
rect 1839 831 2031 837
rect 1839 797 1851 831
rect 2019 797 2031 831
rect 1839 791 2031 797
rect -2087 738 -2041 750
rect -2087 -738 -2081 738
rect -2047 -738 -2041 738
rect -2087 -750 -2041 -738
rect -1829 738 -1783 750
rect -1829 -738 -1823 738
rect -1789 -738 -1783 738
rect -1829 -750 -1783 -738
rect -1571 738 -1525 750
rect -1571 -738 -1565 738
rect -1531 -738 -1525 738
rect -1571 -750 -1525 -738
rect -1313 738 -1267 750
rect -1313 -738 -1307 738
rect -1273 -738 -1267 738
rect -1313 -750 -1267 -738
rect -1055 738 -1009 750
rect -1055 -738 -1049 738
rect -1015 -738 -1009 738
rect -1055 -750 -1009 -738
rect -797 738 -751 750
rect -797 -738 -791 738
rect -757 -738 -751 738
rect -797 -750 -751 -738
rect -539 738 -493 750
rect -539 -738 -533 738
rect -499 -738 -493 738
rect -539 -750 -493 -738
rect -281 738 -235 750
rect -281 -738 -275 738
rect -241 -738 -235 738
rect -281 -750 -235 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 235 738 281 750
rect 235 -738 241 738
rect 275 -738 281 738
rect 235 -750 281 -738
rect 493 738 539 750
rect 493 -738 499 738
rect 533 -738 539 738
rect 493 -750 539 -738
rect 751 738 797 750
rect 751 -738 757 738
rect 791 -738 797 738
rect 751 -750 797 -738
rect 1009 738 1055 750
rect 1009 -738 1015 738
rect 1049 -738 1055 738
rect 1009 -750 1055 -738
rect 1267 738 1313 750
rect 1267 -738 1273 738
rect 1307 -738 1313 738
rect 1267 -750 1313 -738
rect 1525 738 1571 750
rect 1525 -738 1531 738
rect 1565 -738 1571 738
rect 1525 -750 1571 -738
rect 1783 738 1829 750
rect 1783 -738 1789 738
rect 1823 -738 1829 738
rect 1783 -750 1829 -738
rect 2041 738 2087 750
rect 2041 -738 2047 738
rect 2081 -738 2087 738
rect 2041 -750 2087 -738
rect -2031 -797 -1839 -791
rect -2031 -831 -2019 -797
rect -1851 -831 -1839 -797
rect -2031 -837 -1839 -831
rect -1773 -797 -1581 -791
rect -1773 -831 -1761 -797
rect -1593 -831 -1581 -797
rect -1773 -837 -1581 -831
rect -1515 -797 -1323 -791
rect -1515 -831 -1503 -797
rect -1335 -831 -1323 -797
rect -1515 -837 -1323 -831
rect -1257 -797 -1065 -791
rect -1257 -831 -1245 -797
rect -1077 -831 -1065 -797
rect -1257 -837 -1065 -831
rect -999 -797 -807 -791
rect -999 -831 -987 -797
rect -819 -831 -807 -797
rect -999 -837 -807 -831
rect -741 -797 -549 -791
rect -741 -831 -729 -797
rect -561 -831 -549 -797
rect -741 -837 -549 -831
rect -483 -797 -291 -791
rect -483 -831 -471 -797
rect -303 -831 -291 -797
rect -483 -837 -291 -831
rect -225 -797 -33 -791
rect -225 -831 -213 -797
rect -45 -831 -33 -797
rect -225 -837 -33 -831
rect 33 -797 225 -791
rect 33 -831 45 -797
rect 213 -831 225 -797
rect 33 -837 225 -831
rect 291 -797 483 -791
rect 291 -831 303 -797
rect 471 -831 483 -797
rect 291 -837 483 -831
rect 549 -797 741 -791
rect 549 -831 561 -797
rect 729 -831 741 -797
rect 549 -837 741 -831
rect 807 -797 999 -791
rect 807 -831 819 -797
rect 987 -831 999 -797
rect 807 -837 999 -831
rect 1065 -797 1257 -791
rect 1065 -831 1077 -797
rect 1245 -831 1257 -797
rect 1065 -837 1257 -831
rect 1323 -797 1515 -791
rect 1323 -831 1335 -797
rect 1503 -831 1515 -797
rect 1323 -837 1515 -831
rect 1581 -797 1773 -791
rect 1581 -831 1593 -797
rect 1761 -831 1773 -797
rect 1581 -837 1773 -831
rect 1839 -797 2031 -791
rect 1839 -831 1851 -797
rect 2019 -831 2031 -797
rect 1839 -837 2031 -831
<< labels >>
rlabel mvnsubdiffcont 0 -952 0 -952 0 B
port 1 nsew
rlabel mvpdiffc -2064 0 -2064 0 0 D0
port 2 nsew
rlabel polycont -1935 814 -1935 814 0 G0
port 3 nsew
rlabel mvpdiffc -1806 0 -1806 0 0 S1
port 4 nsew
rlabel polycont -1677 814 -1677 814 0 G1
port 5 nsew
rlabel mvpdiffc -1548 0 -1548 0 0 D2
port 6 nsew
rlabel polycont -1419 814 -1419 814 0 G2
port 7 nsew
rlabel mvpdiffc -1290 0 -1290 0 0 S3
port 8 nsew
rlabel polycont -1161 814 -1161 814 0 G3
port 9 nsew
rlabel mvpdiffc -1032 0 -1032 0 0 D4
port 10 nsew
rlabel polycont -903 814 -903 814 0 G4
port 11 nsew
rlabel mvpdiffc -774 0 -774 0 0 S5
port 12 nsew
rlabel polycont -645 814 -645 814 0 G5
port 13 nsew
rlabel mvpdiffc -516 0 -516 0 0 D6
port 14 nsew
rlabel polycont -387 814 -387 814 0 G6
port 15 nsew
rlabel mvpdiffc -258 0 -258 0 0 S7
port 16 nsew
rlabel polycont -129 814 -129 814 0 G7
port 17 nsew
rlabel mvpdiffc 0 0 0 0 0 D8
port 18 nsew
rlabel polycont 129 814 129 814 0 G8
port 19 nsew
rlabel mvpdiffc 258 0 258 0 0 S9
port 20 nsew
rlabel polycont 387 814 387 814 0 G9
port 21 nsew
rlabel mvpdiffc 516 0 516 0 0 D10
port 22 nsew
rlabel polycont 645 814 645 814 0 G10
port 23 nsew
rlabel mvpdiffc 774 0 774 0 0 S11
port 24 nsew
rlabel polycont 903 814 903 814 0 G11
port 25 nsew
rlabel mvpdiffc 1032 0 1032 0 0 D12
port 26 nsew
rlabel polycont 1161 814 1161 814 0 G12
port 27 nsew
rlabel mvpdiffc 1290 0 1290 0 0 S13
port 28 nsew
rlabel polycont 1419 814 1419 814 0 G13
port 29 nsew
rlabel mvpdiffc 1548 0 1548 0 0 D14
port 30 nsew
rlabel polycont 1677 814 1677 814 0 G14
port 31 nsew
rlabel mvpdiffc 1806 0 1806 0 0 S15
port 32 nsew
rlabel polycont 1935 814 1935 814 0 G15
port 33 nsew
<< properties >>
string FIXED_BBOX -2198 -952 2198 952
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
