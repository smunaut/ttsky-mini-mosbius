magic
tech sky130A
magscale 1 2
timestamp 1756580837
<< viali >>
rect 1101 12534 6259 12568
rect 1001 10730 1035 12468
rect 6325 10730 6359 12468
rect 1101 10630 6259 10664
<< metal1 >>
rect 4340 12574 4346 12577
rect 995 12568 4346 12574
rect 4574 12574 4580 12577
rect 4574 12568 6365 12574
rect 995 12534 1101 12568
rect 6259 12534 6365 12568
rect 995 12528 4346 12534
rect 995 12468 1041 12528
rect 4340 12525 4346 12528
rect 4574 12528 6365 12534
rect 4574 12525 4580 12528
rect 995 10730 1001 12468
rect 1035 10730 1041 12468
rect 1205 12485 1257 12491
rect 1363 12485 1415 12491
rect 1277 12390 1343 12436
rect 1837 12485 1889 12491
rect 1593 12390 1659 12436
rect 1995 12485 2047 12491
rect 1521 12335 1573 12341
rect 1909 12390 1975 12436
rect 2469 12485 2521 12491
rect 1679 12335 1731 12341
rect 2225 12390 2291 12436
rect 2627 12485 2679 12491
rect 2153 12335 2205 12341
rect 2541 12390 2607 12436
rect 3101 12485 3153 12491
rect 2311 12335 2363 12341
rect 2857 12390 2923 12436
rect 3259 12485 3311 12491
rect 2785 12335 2837 12341
rect 3173 12390 3239 12436
rect 4049 12485 4101 12491
rect 2943 12335 2995 12341
rect 3489 12390 3555 12436
rect 3417 12335 3469 12341
rect 3575 12335 3627 12341
rect 3805 12390 3871 12436
rect 4207 12485 4259 12491
rect 3733 12335 3785 12341
rect 4121 12390 4187 12436
rect 4681 12485 4733 12491
rect 3891 12335 3943 12341
rect 4437 12390 4503 12436
rect 4839 12485 4891 12491
rect 4365 12335 4417 12341
rect 4753 12390 4819 12436
rect 5313 12485 5365 12491
rect 4523 12335 4575 12341
rect 5069 12390 5135 12436
rect 5471 12485 5523 12491
rect 4997 12335 5049 12341
rect 5385 12390 5451 12436
rect 5945 12485 5997 12491
rect 5155 12335 5207 12341
rect 5701 12390 5767 12436
rect 6103 12485 6155 12491
rect 5629 12335 5681 12341
rect 6017 12390 6083 12436
rect 6319 12468 6365 12528
rect 5787 12335 5839 12341
rect 1126 12043 1178 12049
rect 1126 11149 1178 11155
rect 1284 12043 1336 12049
rect 1284 11149 1336 11155
rect 1442 12043 1494 12049
rect 1442 11149 1494 11155
rect 1600 12043 1652 12049
rect 1600 11149 1652 11155
rect 1758 12043 1810 12049
rect 1758 11149 1810 11155
rect 1916 12043 1968 12049
rect 1916 11149 1968 11155
rect 2074 12043 2126 12049
rect 2074 11149 2126 11155
rect 2232 12043 2284 12049
rect 2232 11149 2284 11155
rect 2390 12043 2442 12049
rect 2390 11149 2442 11155
rect 2548 12043 2600 12049
rect 2548 11149 2600 11155
rect 2706 12043 2758 12049
rect 2706 11149 2758 11155
rect 2864 12043 2916 12049
rect 2864 11149 2916 11155
rect 3022 12043 3074 12049
rect 3022 11149 3074 11155
rect 3180 12043 3232 12049
rect 3180 11149 3232 11155
rect 3338 12043 3390 12049
rect 3338 11149 3390 11155
rect 3496 12043 3548 12049
rect 3496 11149 3548 11155
rect 3654 12043 3706 12049
rect 3654 11149 3706 11155
rect 3812 12043 3864 12049
rect 3812 11149 3864 11155
rect 3970 12043 4022 12049
rect 3970 11149 4022 11155
rect 4128 12043 4180 12049
rect 4128 11149 4180 11155
rect 4286 12043 4338 12049
rect 4286 11149 4338 11155
rect 4444 12043 4496 12049
rect 4444 11149 4496 11155
rect 4602 12043 4654 12049
rect 4602 11149 4654 11155
rect 4760 12043 4812 12049
rect 4760 11149 4812 11155
rect 4918 12043 4970 12049
rect 4918 11149 4970 11155
rect 5076 12043 5128 12049
rect 5076 11149 5128 11155
rect 5234 12043 5286 12049
rect 5234 11149 5286 11155
rect 5392 12043 5444 12049
rect 5392 11149 5444 11155
rect 5550 12043 5602 12049
rect 5550 11149 5602 11155
rect 5708 12043 5760 12049
rect 5708 11149 5760 11155
rect 5866 12043 5918 12049
rect 5866 11149 5918 11155
rect 6024 12043 6076 12049
rect 6024 11149 6076 11155
rect 6182 12043 6234 12049
rect 6182 11149 6234 11155
rect 1205 10857 1257 10863
rect 1363 10857 1415 10863
rect 1277 10762 1343 10808
rect 1837 10857 1889 10863
rect 995 10670 1041 10730
rect 1593 10762 1659 10808
rect 1995 10857 2047 10863
rect 1521 10707 1573 10713
rect 1909 10762 1975 10808
rect 2469 10857 2521 10863
rect 1679 10707 1731 10713
rect 2225 10762 2291 10808
rect 2627 10857 2679 10863
rect 2153 10707 2205 10713
rect 2541 10762 2607 10808
rect 3101 10857 3153 10863
rect 2311 10707 2363 10713
rect 2857 10762 2923 10808
rect 3259 10857 3311 10863
rect 2785 10707 2837 10713
rect 3173 10762 3239 10808
rect 4049 10857 4101 10863
rect 2943 10707 2995 10713
rect 3489 10762 3555 10808
rect 3417 10707 3469 10713
rect 3575 10707 3627 10713
rect 3805 10762 3871 10808
rect 4207 10857 4259 10863
rect 3733 10707 3785 10713
rect 4121 10762 4187 10808
rect 4681 10857 4733 10863
rect 3891 10707 3943 10713
rect 4437 10762 4503 10808
rect 4839 10857 4891 10863
rect 4365 10707 4417 10713
rect 4753 10762 4819 10808
rect 5313 10857 5365 10863
rect 4523 10707 4575 10713
rect 5069 10762 5135 10808
rect 5471 10857 5523 10863
rect 4997 10707 5049 10713
rect 5385 10762 5451 10808
rect 5945 10857 5997 10863
rect 5155 10707 5207 10713
rect 5701 10762 5767 10808
rect 6103 10857 6155 10863
rect 5629 10707 5681 10713
rect 6017 10762 6083 10808
rect 5787 10707 5839 10713
rect 6319 10730 6325 12468
rect 6359 10730 6365 12468
rect 4340 10670 4346 10673
rect 995 10664 4346 10670
rect 4574 10670 4580 10673
rect 6319 10670 6365 10730
rect 4574 10664 6365 10670
rect 995 10630 1101 10664
rect 6259 10630 6365 10664
rect 995 10624 4346 10630
rect 4340 10621 4346 10624
rect 4574 10624 6365 10630
rect 4574 10621 4580 10624
<< via1 >>
rect 4346 12568 4574 12577
rect 4346 12534 4574 12568
rect 4346 12525 4574 12534
rect 1205 12433 1257 12485
rect 1363 12433 1415 12485
rect 1521 12341 1573 12393
rect 1837 12433 1889 12485
rect 1679 12341 1731 12393
rect 1995 12433 2047 12485
rect 2153 12341 2205 12393
rect 2469 12433 2521 12485
rect 2311 12341 2363 12393
rect 2627 12433 2679 12485
rect 2785 12341 2837 12393
rect 3101 12433 3153 12485
rect 2943 12341 2995 12393
rect 3259 12433 3311 12485
rect 3417 12341 3469 12393
rect 3575 12341 3627 12393
rect 3733 12341 3785 12393
rect 4049 12433 4101 12485
rect 3891 12341 3943 12393
rect 4207 12433 4259 12485
rect 4365 12341 4417 12393
rect 4681 12433 4733 12485
rect 4523 12341 4575 12393
rect 4839 12433 4891 12485
rect 4997 12341 5049 12393
rect 5313 12433 5365 12485
rect 5155 12341 5207 12393
rect 5471 12433 5523 12485
rect 5629 12341 5681 12393
rect 5945 12433 5997 12485
rect 5787 12341 5839 12393
rect 6103 12433 6155 12485
rect 1126 11155 1178 12043
rect 1284 11155 1336 12043
rect 1442 11155 1494 12043
rect 1600 11155 1652 12043
rect 1758 11155 1810 12043
rect 1916 11155 1968 12043
rect 2074 11155 2126 12043
rect 2232 11155 2284 12043
rect 2390 11155 2442 12043
rect 2548 11155 2600 12043
rect 2706 11155 2758 12043
rect 2864 11155 2916 12043
rect 3022 11155 3074 12043
rect 3180 11155 3232 12043
rect 3338 11155 3390 12043
rect 3496 11155 3548 12043
rect 3654 11155 3706 12043
rect 3812 11155 3864 12043
rect 3970 11155 4022 12043
rect 4128 11155 4180 12043
rect 4286 11155 4338 12043
rect 4444 11155 4496 12043
rect 4602 11155 4654 12043
rect 4760 11155 4812 12043
rect 4918 11155 4970 12043
rect 5076 11155 5128 12043
rect 5234 11155 5286 12043
rect 5392 11155 5444 12043
rect 5550 11155 5602 12043
rect 5708 11155 5760 12043
rect 5866 11155 5918 12043
rect 6024 11155 6076 12043
rect 6182 11155 6234 12043
rect 1205 10805 1257 10857
rect 1363 10805 1415 10857
rect 1521 10713 1573 10765
rect 1837 10805 1889 10857
rect 1679 10713 1731 10765
rect 1995 10805 2047 10857
rect 2153 10713 2205 10765
rect 2469 10805 2521 10857
rect 2311 10713 2363 10765
rect 2627 10805 2679 10857
rect 2785 10713 2837 10765
rect 3101 10805 3153 10857
rect 2943 10713 2995 10765
rect 3259 10805 3311 10857
rect 3417 10713 3469 10765
rect 3575 10713 3627 10765
rect 3733 10713 3785 10765
rect 4049 10805 4101 10857
rect 3891 10713 3943 10765
rect 4207 10805 4259 10857
rect 4365 10713 4417 10765
rect 4681 10805 4733 10857
rect 4523 10713 4575 10765
rect 4839 10805 4891 10857
rect 4997 10713 5049 10765
rect 5313 10805 5365 10857
rect 5155 10713 5207 10765
rect 5471 10805 5523 10857
rect 5629 10713 5681 10765
rect 5945 10805 5997 10857
rect 5787 10713 5839 10765
rect 6103 10805 6155 10857
rect 4346 10664 4574 10673
rect 4346 10630 4574 10664
rect 4346 10621 4574 10630
<< metal2 >>
rect 992 12691 1128 12700
rect 6232 12599 6368 12608
rect 4340 12577 4349 12579
rect 4571 12577 4580 12579
rect 4340 12525 4346 12577
rect 4574 12525 4580 12577
rect 4340 12523 4349 12525
rect 4571 12523 4580 12525
rect 992 12485 1128 12501
rect 992 12433 1205 12485
rect 1257 12433 1363 12485
rect 1415 12433 1837 12485
rect 1889 12433 1995 12485
rect 2047 12433 2469 12485
rect 2521 12433 2627 12485
rect 2679 12433 3101 12485
rect 3153 12433 3259 12485
rect 3311 12433 4049 12485
rect 4101 12433 4207 12485
rect 4259 12433 4681 12485
rect 4733 12433 4839 12485
rect 4891 12433 5313 12485
rect 5365 12433 5471 12485
rect 5523 12433 5945 12485
rect 5997 12433 6103 12485
rect 6155 12433 6175 12485
rect 992 10857 1044 12433
rect 6232 12393 6368 12409
rect 1185 12341 1521 12393
rect 1573 12341 1679 12393
rect 1731 12341 2153 12393
rect 2205 12341 2311 12393
rect 2363 12341 2785 12393
rect 2837 12341 2943 12393
rect 2995 12341 3417 12393
rect 3469 12341 3575 12393
rect 3627 12341 3733 12393
rect 3785 12341 3891 12393
rect 3943 12341 4365 12393
rect 4417 12341 4523 12393
rect 4575 12341 4997 12393
rect 5049 12341 5155 12393
rect 5207 12341 5629 12393
rect 5681 12341 5787 12393
rect 5839 12341 6368 12393
rect 1126 12043 1178 12049
rect 1124 11744 1126 11753
rect 1284 12043 1336 12049
rect 1178 11744 1180 11753
rect 1124 11445 1126 11454
rect 1178 11445 1180 11454
rect 1126 11149 1178 11155
rect 1244 11344 1284 11353
rect 1442 12043 1494 12049
rect 1400 11744 1442 11753
rect 1560 12044 1696 12053
rect 1560 11845 1600 11854
rect 1494 11744 1536 11753
rect 1400 11445 1442 11454
rect 1336 11344 1380 11353
rect 1244 11145 1380 11154
rect 1494 11445 1536 11454
rect 1442 11149 1494 11155
rect 1652 11845 1696 11854
rect 1758 12043 1810 12049
rect 1716 11744 1758 11753
rect 1916 12043 1968 12049
rect 1810 11744 1852 11753
rect 1716 11445 1758 11454
rect 1600 11149 1652 11155
rect 1810 11445 1852 11454
rect 1758 11149 1810 11155
rect 1876 11344 1916 11353
rect 2074 12043 2126 12049
rect 2032 11744 2074 11753
rect 2192 12044 2328 12053
rect 2192 11845 2232 11854
rect 2126 11744 2168 11753
rect 2032 11445 2074 11454
rect 1968 11344 2012 11353
rect 1876 11145 2012 11154
rect 2126 11445 2168 11454
rect 2074 11149 2126 11155
rect 2284 11845 2328 11854
rect 2390 12043 2442 12049
rect 2348 11744 2390 11753
rect 2548 12043 2600 12049
rect 2442 11744 2484 11753
rect 2348 11445 2390 11454
rect 2232 11149 2284 11155
rect 2442 11445 2484 11454
rect 2390 11149 2442 11155
rect 2508 11344 2548 11353
rect 2706 12043 2758 12049
rect 2664 11744 2706 11753
rect 2824 12044 2960 12053
rect 2824 11845 2864 11854
rect 2758 11744 2800 11753
rect 2664 11445 2706 11454
rect 2600 11344 2644 11353
rect 2508 11145 2644 11154
rect 2758 11445 2800 11454
rect 2706 11149 2758 11155
rect 2916 11845 2960 11854
rect 3022 12043 3074 12049
rect 2980 11744 3022 11753
rect 3180 12043 3232 12049
rect 3074 11744 3116 11753
rect 2980 11445 3022 11454
rect 2864 11149 2916 11155
rect 3074 11445 3116 11454
rect 3022 11149 3074 11155
rect 3140 11344 3180 11353
rect 3338 12043 3390 12049
rect 3296 11744 3338 11753
rect 3456 12044 3592 12053
rect 3456 11845 3496 11854
rect 3390 11744 3432 11753
rect 3296 11445 3338 11454
rect 3232 11344 3276 11353
rect 3140 11145 3276 11154
rect 3390 11445 3432 11454
rect 3338 11149 3390 11155
rect 3548 11845 3592 11854
rect 3654 12043 3706 12049
rect 3612 11744 3654 11753
rect 3772 12044 3908 12053
rect 3772 11845 3812 11854
rect 3706 11744 3748 11753
rect 3612 11445 3654 11454
rect 3496 11149 3548 11155
rect 3706 11445 3748 11454
rect 3654 11149 3706 11155
rect 3864 11845 3908 11854
rect 3970 12043 4022 12049
rect 3928 11744 3970 11753
rect 4128 12043 4180 12049
rect 4022 11744 4064 11753
rect 3928 11445 3970 11454
rect 3812 11149 3864 11155
rect 4022 11445 4064 11454
rect 3970 11149 4022 11155
rect 4088 11344 4128 11353
rect 4286 12043 4338 12049
rect 4244 11744 4286 11753
rect 4404 12044 4540 12053
rect 4404 11845 4444 11854
rect 4338 11744 4380 11753
rect 4244 11445 4286 11454
rect 4180 11344 4224 11353
rect 4088 11145 4224 11154
rect 4338 11445 4380 11454
rect 4286 11149 4338 11155
rect 4496 11845 4540 11854
rect 4602 12043 4654 12049
rect 4560 11744 4602 11753
rect 4760 12043 4812 12049
rect 4654 11744 4696 11753
rect 4560 11445 4602 11454
rect 4444 11149 4496 11155
rect 4654 11445 4696 11454
rect 4602 11149 4654 11155
rect 4720 11344 4760 11353
rect 4918 12043 4970 12049
rect 4876 11744 4918 11753
rect 5036 12044 5172 12053
rect 5036 11845 5076 11854
rect 4970 11744 5012 11753
rect 4876 11445 4918 11454
rect 4812 11344 4856 11353
rect 4720 11145 4856 11154
rect 4970 11445 5012 11454
rect 4918 11149 4970 11155
rect 5128 11845 5172 11854
rect 5234 12043 5286 12049
rect 5192 11744 5234 11753
rect 5392 12043 5444 12049
rect 5286 11744 5328 11753
rect 5192 11445 5234 11454
rect 5076 11149 5128 11155
rect 5286 11445 5328 11454
rect 5234 11149 5286 11155
rect 5352 11344 5392 11353
rect 5550 12043 5602 12049
rect 5508 11744 5550 11753
rect 5668 12044 5804 12053
rect 5668 11845 5708 11854
rect 5602 11744 5644 11753
rect 5508 11445 5550 11454
rect 5444 11344 5488 11353
rect 5352 11145 5488 11154
rect 5602 11445 5644 11454
rect 5550 11149 5602 11155
rect 5760 11845 5804 11854
rect 5866 12043 5918 12049
rect 5824 11744 5866 11753
rect 6024 12043 6076 12049
rect 5918 11744 5960 11753
rect 5824 11445 5866 11454
rect 5708 11149 5760 11155
rect 5918 11445 5960 11454
rect 5866 11149 5918 11155
rect 5984 11344 6024 11353
rect 6182 12043 6234 12049
rect 6180 11744 6182 11753
rect 6234 11744 6236 11753
rect 6180 11445 6182 11454
rect 6076 11344 6120 11353
rect 5984 11145 6120 11154
rect 6234 11445 6236 11454
rect 6182 11149 6234 11155
rect 992 10805 1205 10857
rect 1257 10805 1363 10857
rect 1415 10805 1837 10857
rect 1889 10805 1995 10857
rect 2047 10805 2469 10857
rect 2521 10805 2627 10857
rect 2679 10805 3101 10857
rect 3153 10805 3259 10857
rect 3311 10805 4049 10857
rect 4101 10805 4207 10857
rect 4259 10805 4681 10857
rect 4733 10805 4839 10857
rect 4891 10805 5313 10857
rect 5365 10805 5471 10857
rect 5523 10805 5945 10857
rect 5997 10805 6103 10857
rect 6155 10805 6175 10857
rect 6316 10765 6368 12341
rect 1185 10713 1521 10765
rect 1573 10713 1679 10765
rect 1731 10713 2153 10765
rect 2205 10713 2311 10765
rect 2363 10713 2785 10765
rect 2837 10713 2943 10765
rect 2995 10713 3417 10765
rect 3469 10713 3575 10765
rect 3627 10713 3733 10765
rect 3785 10713 3891 10765
rect 3943 10713 4365 10765
rect 4417 10713 4523 10765
rect 4575 10713 4997 10765
rect 5049 10713 5155 10765
rect 5207 10713 5629 10765
rect 5681 10713 5787 10765
rect 5839 10713 6368 10765
rect 4340 10673 4349 10675
rect 4571 10673 4580 10675
rect 4340 10621 4346 10673
rect 4574 10621 4580 10673
rect 4340 10619 4349 10621
rect 4571 10619 4580 10621
<< via2 >>
rect 992 12501 1128 12691
rect 4349 12577 4571 12579
rect 4349 12525 4571 12577
rect 4349 12523 4571 12525
rect 6232 12409 6368 12599
rect 1124 11454 1126 11744
rect 1126 11454 1178 11744
rect 1178 11454 1180 11744
rect 1560 12043 1696 12044
rect 1560 11854 1600 12043
rect 1600 11854 1652 12043
rect 1652 11854 1696 12043
rect 1400 11454 1442 11744
rect 1442 11454 1494 11744
rect 1494 11454 1536 11744
rect 1244 11155 1284 11344
rect 1284 11155 1336 11344
rect 1336 11155 1380 11344
rect 1244 11154 1380 11155
rect 1716 11454 1758 11744
rect 1758 11454 1810 11744
rect 1810 11454 1852 11744
rect 2192 12043 2328 12044
rect 2192 11854 2232 12043
rect 2232 11854 2284 12043
rect 2284 11854 2328 12043
rect 2032 11454 2074 11744
rect 2074 11454 2126 11744
rect 2126 11454 2168 11744
rect 1876 11155 1916 11344
rect 1916 11155 1968 11344
rect 1968 11155 2012 11344
rect 1876 11154 2012 11155
rect 2348 11454 2390 11744
rect 2390 11454 2442 11744
rect 2442 11454 2484 11744
rect 2824 12043 2960 12044
rect 2824 11854 2864 12043
rect 2864 11854 2916 12043
rect 2916 11854 2960 12043
rect 2664 11454 2706 11744
rect 2706 11454 2758 11744
rect 2758 11454 2800 11744
rect 2508 11155 2548 11344
rect 2548 11155 2600 11344
rect 2600 11155 2644 11344
rect 2508 11154 2644 11155
rect 2980 11454 3022 11744
rect 3022 11454 3074 11744
rect 3074 11454 3116 11744
rect 3456 12043 3592 12044
rect 3456 11854 3496 12043
rect 3496 11854 3548 12043
rect 3548 11854 3592 12043
rect 3296 11454 3338 11744
rect 3338 11454 3390 11744
rect 3390 11454 3432 11744
rect 3140 11155 3180 11344
rect 3180 11155 3232 11344
rect 3232 11155 3276 11344
rect 3140 11154 3276 11155
rect 3772 12043 3908 12044
rect 3772 11854 3812 12043
rect 3812 11854 3864 12043
rect 3864 11854 3908 12043
rect 3612 11454 3654 11744
rect 3654 11454 3706 11744
rect 3706 11454 3748 11744
rect 3928 11454 3970 11744
rect 3970 11454 4022 11744
rect 4022 11454 4064 11744
rect 4404 12043 4540 12044
rect 4404 11854 4444 12043
rect 4444 11854 4496 12043
rect 4496 11854 4540 12043
rect 4244 11454 4286 11744
rect 4286 11454 4338 11744
rect 4338 11454 4380 11744
rect 4088 11155 4128 11344
rect 4128 11155 4180 11344
rect 4180 11155 4224 11344
rect 4088 11154 4224 11155
rect 4560 11454 4602 11744
rect 4602 11454 4654 11744
rect 4654 11454 4696 11744
rect 5036 12043 5172 12044
rect 5036 11854 5076 12043
rect 5076 11854 5128 12043
rect 5128 11854 5172 12043
rect 4876 11454 4918 11744
rect 4918 11454 4970 11744
rect 4970 11454 5012 11744
rect 4720 11155 4760 11344
rect 4760 11155 4812 11344
rect 4812 11155 4856 11344
rect 4720 11154 4856 11155
rect 5192 11454 5234 11744
rect 5234 11454 5286 11744
rect 5286 11454 5328 11744
rect 5668 12043 5804 12044
rect 5668 11854 5708 12043
rect 5708 11854 5760 12043
rect 5760 11854 5804 12043
rect 5508 11454 5550 11744
rect 5550 11454 5602 11744
rect 5602 11454 5644 11744
rect 5352 11155 5392 11344
rect 5392 11155 5444 11344
rect 5444 11155 5488 11344
rect 5352 11154 5488 11155
rect 5824 11454 5866 11744
rect 5866 11454 5918 11744
rect 5918 11454 5960 11744
rect 6180 11454 6182 11744
rect 6182 11454 6234 11744
rect 6234 11454 6236 11744
rect 5984 11155 6024 11344
rect 6024 11155 6076 11344
rect 6076 11155 6120 11344
rect 5984 11154 6120 11155
rect 4349 10673 4571 10675
rect 4349 10621 4571 10673
rect 4349 10619 4571 10621
<< metal3 >>
rect 987 12843 2590 12844
rect 987 12699 2296 12843
rect 2584 12699 2590 12843
rect 987 12698 2590 12699
rect 2890 12843 6373 12844
rect 2890 12699 2896 12843
rect 3184 12699 6373 12843
rect 2890 12698 6373 12699
rect 987 12691 1133 12698
rect 987 12501 992 12691
rect 1128 12501 1133 12691
rect 6227 12599 6373 12698
rect 4340 12583 4580 12584
rect 4340 12519 4346 12583
rect 4574 12519 4580 12583
rect 4340 12518 4580 12519
rect 987 12496 1133 12501
rect 6227 12409 6232 12599
rect 6368 12409 6373 12599
rect 6227 12404 6373 12409
rect 1555 12044 7170 12049
rect 1555 11854 1560 12044
rect 1696 11854 2192 12044
rect 2328 11854 2824 12044
rect 2960 11854 3456 12044
rect 3592 11854 3772 12044
rect 3908 11854 4404 12044
rect 4540 11854 5036 12044
rect 5172 11854 5668 12044
rect 5804 11854 7170 12044
rect 1555 11849 7170 11854
rect 1119 11748 6241 11749
rect 1119 11744 2891 11748
rect 3189 11744 6241 11748
rect 1119 11454 1124 11744
rect 1180 11454 1400 11744
rect 1536 11454 1716 11744
rect 1852 11454 2032 11744
rect 2168 11454 2348 11744
rect 2484 11454 2664 11744
rect 2800 11454 2891 11744
rect 3189 11454 3296 11744
rect 3432 11454 3612 11744
rect 3748 11454 3928 11744
rect 4064 11454 4244 11744
rect 4380 11454 4560 11744
rect 4696 11454 4876 11744
rect 5012 11454 5192 11744
rect 5328 11454 5508 11744
rect 5644 11454 5824 11744
rect 5960 11454 6180 11744
rect 6236 11454 6241 11744
rect 1119 11450 2891 11454
rect 3189 11450 6241 11454
rect 1119 11449 6241 11450
rect 1239 11348 6270 11349
rect 1239 11344 5976 11348
rect 1239 11154 1244 11344
rect 1380 11154 1876 11344
rect 2012 11154 2508 11344
rect 2644 11154 3140 11344
rect 3276 11154 4088 11344
rect 4224 11154 4720 11344
rect 4856 11154 5352 11344
rect 5488 11154 5976 11344
rect 1239 11150 5976 11154
rect 6264 11150 6270 11348
rect 1239 11149 6270 11150
rect 4340 10679 4580 10680
rect 4340 10615 4346 10679
rect 4574 10615 4580 10679
rect 4340 10614 4580 10615
rect 6970 10114 7170 11849
rect 6970 10113 9950 10114
rect 6970 9915 9656 10113
rect 9944 9915 9950 10113
rect 6970 9914 9950 9915
rect 7292 8249 10550 8250
rect 7292 7851 10256 8249
rect 10544 7851 10550 8249
rect 7292 7850 10550 7851
rect 954 5846 1001 5910
rect 1065 5846 1071 5910
rect 4634 5846 4681 5910
rect 4745 5846 4751 5910
rect 954 1224 1121 1288
rect 1185 1224 1191 1288
rect 4634 1224 4801 1288
rect 4865 1224 4871 1288
<< via3 >>
rect 2296 12699 2584 12843
rect 2896 12699 3184 12843
rect 4346 12579 4574 12583
rect 4346 12523 4349 12579
rect 4349 12523 4571 12579
rect 4571 12523 4574 12579
rect 4346 12519 4574 12523
rect 2891 11744 3189 11748
rect 2891 11454 2980 11744
rect 2980 11454 3116 11744
rect 3116 11454 3189 11744
rect 2891 11450 3189 11454
rect 5976 11344 6264 11348
rect 5976 11154 5984 11344
rect 5984 11154 6120 11344
rect 6120 11154 6264 11344
rect 5976 11150 6264 11154
rect 4346 10675 4574 10679
rect 4346 10619 4349 10675
rect 4349 10619 4571 10675
rect 4571 10619 4574 10675
rect 4346 10615 4574 10619
rect 9656 9915 9944 10113
rect 661 7851 899 8249
rect 4341 7851 4579 8249
rect 10256 7851 10544 8249
rect 2891 6147 3189 6545
rect 1001 5846 1065 5910
rect 4681 5846 4745 5910
rect 661 3229 899 3627
rect 4341 3229 4579 3627
rect 2291 1525 2589 1923
rect 6571 1525 6869 1923
rect 1121 1224 1185 1288
rect 4801 1224 4865 1288
<< metal4 >>
rect 20 10198 260 12998
rect 340 10198 580 12998
rect 660 10198 900 12998
rect 1690 9200 1990 12998
rect 2290 12843 2590 12998
rect 2290 12699 2296 12843
rect 2584 12699 2590 12843
rect 2290 12698 2590 12699
rect 2890 12843 3190 12998
rect 2890 12699 2896 12843
rect 3184 12699 3190 12843
rect 2890 12698 3190 12699
rect 2890 11748 3190 11749
rect 2890 11450 2891 11748
rect 3189 11450 3190 11748
rect 1690 8900 2590 9200
rect 1000 5910 1066 5911
rect 1000 5846 1001 5910
rect 1065 5846 1066 5910
rect 20 5576 260 5846
rect 340 5576 580 5846
rect 660 5576 900 5846
rect 1000 5845 1066 5846
rect 20 1136 260 1224
rect 340 1136 580 1224
rect 660 -48 900 1224
rect 1000 1140 1060 5845
rect 2290 1923 2590 8900
rect 2890 6545 3190 11450
rect 3700 10198 3940 12998
rect 4020 10198 4260 12998
rect 4340 12583 4580 12998
rect 4340 12519 4346 12583
rect 4574 12519 4580 12583
rect 4340 10679 4580 12519
rect 5970 11348 6270 12998
rect 5970 11150 5976 11348
rect 6264 11150 6270 11348
rect 5970 11149 6270 11150
rect 4340 10615 4346 10679
rect 4574 10615 4580 10679
rect 4340 10198 4580 10615
rect 2890 6147 2891 6545
rect 3189 6147 3190 6545
rect 2890 6146 3190 6147
rect 4680 5910 4746 5911
rect 4680 5846 4681 5910
rect 4745 5846 4746 5910
rect 3700 5576 3940 5846
rect 4020 5576 4260 5846
rect 4340 5576 4580 5846
rect 4680 5845 4746 5846
rect 2290 1525 2291 1923
rect 2589 1525 2590 1923
rect 2290 1524 2590 1525
rect 1120 1288 1186 1289
rect 1120 1224 1121 1288
rect 1185 1224 1186 1288
rect 1120 1221 1186 1224
rect 1120 1140 1180 1221
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1140 4740 5845
rect 6570 1923 6870 12998
rect 9650 10113 9950 12998
rect 9650 9915 9656 10113
rect 9944 9915 9950 10113
rect 9650 9914 9950 9915
rect 10250 8249 10550 12998
rect 10250 7851 10256 8249
rect 10544 7851 10550 8249
rect 10250 7850 10550 7851
rect 6570 1525 6571 1923
rect 6869 1525 6870 1923
rect 6570 1524 6870 1525
rect 4800 1288 4866 1289
rect 4800 1224 4801 1288
rect 4865 1224 4866 1288
rect 4800 1221 4866 1224
rect 4800 1140 4860 1221
use dev_ctrl_b2  dev_ctrl_b2_0
timestamp 1756064790
transform 1 0 3680 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e2  dev_ctrl_e2_0
timestamp 1756064830
transform 1 0 0 0 1 0
box -38 -48 6868 1140
use sky130_fd_pr__pfet_g5v0d10v5_GFVKBM  sky130_fd_pr__pfet_g5v0d10v5_GFVKBM_0
timestamp 1756220169
transform 1 0 3680 0 1 11599
box -2757 -1047 2757 1047
use tt_asw_3v3  tt_asw_3v3_0
array 0 1 3680 0 1 -4622
timestamp 1756064685
transform 1 0 0 0 -1 5576
box 0 0 3680 4352
<< end >>
