magic
tech sky130A
magscale 1 2
timestamp 1756064685
<< pwell >>
rect -6909 -758 6909 758
<< mvnmos >>
rect -6679 -500 -6479 500
rect -6421 -500 -6221 500
rect -6163 -500 -5963 500
rect -5905 -500 -5705 500
rect -5647 -500 -5447 500
rect -5389 -500 -5189 500
rect -5131 -500 -4931 500
rect -4873 -500 -4673 500
rect -4615 -500 -4415 500
rect -4357 -500 -4157 500
rect -4099 -500 -3899 500
rect -3841 -500 -3641 500
rect -3583 -500 -3383 500
rect -3325 -500 -3125 500
rect -3067 -500 -2867 500
rect -2809 -500 -2609 500
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
rect 2609 -500 2809 500
rect 2867 -500 3067 500
rect 3125 -500 3325 500
rect 3383 -500 3583 500
rect 3641 -500 3841 500
rect 3899 -500 4099 500
rect 4157 -500 4357 500
rect 4415 -500 4615 500
rect 4673 -500 4873 500
rect 4931 -500 5131 500
rect 5189 -500 5389 500
rect 5447 -500 5647 500
rect 5705 -500 5905 500
rect 5963 -500 6163 500
rect 6221 -500 6421 500
rect 6479 -500 6679 500
<< mvndiff >>
rect -6737 488 -6679 500
rect -6737 -488 -6725 488
rect -6691 -488 -6679 488
rect -6737 -500 -6679 -488
rect -6479 488 -6421 500
rect -6479 -488 -6467 488
rect -6433 -488 -6421 488
rect -6479 -500 -6421 -488
rect -6221 488 -6163 500
rect -6221 -488 -6209 488
rect -6175 -488 -6163 488
rect -6221 -500 -6163 -488
rect -5963 488 -5905 500
rect -5963 -488 -5951 488
rect -5917 -488 -5905 488
rect -5963 -500 -5905 -488
rect -5705 488 -5647 500
rect -5705 -488 -5693 488
rect -5659 -488 -5647 488
rect -5705 -500 -5647 -488
rect -5447 488 -5389 500
rect -5447 -488 -5435 488
rect -5401 -488 -5389 488
rect -5447 -500 -5389 -488
rect -5189 488 -5131 500
rect -5189 -488 -5177 488
rect -5143 -488 -5131 488
rect -5189 -500 -5131 -488
rect -4931 488 -4873 500
rect -4931 -488 -4919 488
rect -4885 -488 -4873 488
rect -4931 -500 -4873 -488
rect -4673 488 -4615 500
rect -4673 -488 -4661 488
rect -4627 -488 -4615 488
rect -4673 -500 -4615 -488
rect -4415 488 -4357 500
rect -4415 -488 -4403 488
rect -4369 -488 -4357 488
rect -4415 -500 -4357 -488
rect -4157 488 -4099 500
rect -4157 -488 -4145 488
rect -4111 -488 -4099 488
rect -4157 -500 -4099 -488
rect -3899 488 -3841 500
rect -3899 -488 -3887 488
rect -3853 -488 -3841 488
rect -3899 -500 -3841 -488
rect -3641 488 -3583 500
rect -3641 -488 -3629 488
rect -3595 -488 -3583 488
rect -3641 -500 -3583 -488
rect -3383 488 -3325 500
rect -3383 -488 -3371 488
rect -3337 -488 -3325 488
rect -3383 -500 -3325 -488
rect -3125 488 -3067 500
rect -3125 -488 -3113 488
rect -3079 -488 -3067 488
rect -3125 -500 -3067 -488
rect -2867 488 -2809 500
rect -2867 -488 -2855 488
rect -2821 -488 -2809 488
rect -2867 -500 -2809 -488
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
rect 2809 488 2867 500
rect 2809 -488 2821 488
rect 2855 -488 2867 488
rect 2809 -500 2867 -488
rect 3067 488 3125 500
rect 3067 -488 3079 488
rect 3113 -488 3125 488
rect 3067 -500 3125 -488
rect 3325 488 3383 500
rect 3325 -488 3337 488
rect 3371 -488 3383 488
rect 3325 -500 3383 -488
rect 3583 488 3641 500
rect 3583 -488 3595 488
rect 3629 -488 3641 488
rect 3583 -500 3641 -488
rect 3841 488 3899 500
rect 3841 -488 3853 488
rect 3887 -488 3899 488
rect 3841 -500 3899 -488
rect 4099 488 4157 500
rect 4099 -488 4111 488
rect 4145 -488 4157 488
rect 4099 -500 4157 -488
rect 4357 488 4415 500
rect 4357 -488 4369 488
rect 4403 -488 4415 488
rect 4357 -500 4415 -488
rect 4615 488 4673 500
rect 4615 -488 4627 488
rect 4661 -488 4673 488
rect 4615 -500 4673 -488
rect 4873 488 4931 500
rect 4873 -488 4885 488
rect 4919 -488 4931 488
rect 4873 -500 4931 -488
rect 5131 488 5189 500
rect 5131 -488 5143 488
rect 5177 -488 5189 488
rect 5131 -500 5189 -488
rect 5389 488 5447 500
rect 5389 -488 5401 488
rect 5435 -488 5447 488
rect 5389 -500 5447 -488
rect 5647 488 5705 500
rect 5647 -488 5659 488
rect 5693 -488 5705 488
rect 5647 -500 5705 -488
rect 5905 488 5963 500
rect 5905 -488 5917 488
rect 5951 -488 5963 488
rect 5905 -500 5963 -488
rect 6163 488 6221 500
rect 6163 -488 6175 488
rect 6209 -488 6221 488
rect 6163 -500 6221 -488
rect 6421 488 6479 500
rect 6421 -488 6433 488
rect 6467 -488 6479 488
rect 6421 -500 6479 -488
rect 6679 488 6737 500
rect 6679 -488 6691 488
rect 6725 -488 6737 488
rect 6679 -500 6737 -488
<< mvndiffc >>
rect -6725 -488 -6691 488
rect -6467 -488 -6433 488
rect -6209 -488 -6175 488
rect -5951 -488 -5917 488
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect 5917 -488 5951 488
rect 6175 -488 6209 488
rect 6433 -488 6467 488
rect 6691 -488 6725 488
<< mvpsubdiff >>
rect -6873 710 6873 722
rect -6873 676 -6765 710
rect 6765 676 6873 710
rect -6873 664 6873 676
rect -6873 614 -6815 664
rect -6873 -614 -6861 614
rect -6827 -614 -6815 614
rect 6815 614 6873 664
rect -6873 -664 -6815 -614
rect 6815 -614 6827 614
rect 6861 -614 6873 614
rect 6815 -664 6873 -614
rect -6873 -676 6873 -664
rect -6873 -710 -6765 -676
rect 6765 -710 6873 -676
rect -6873 -722 6873 -710
<< mvpsubdiffcont >>
rect -6765 676 6765 710
rect -6861 -614 -6827 614
rect 6827 -614 6861 614
rect -6765 -710 6765 -676
<< poly >>
rect -6679 572 -6479 588
rect -6679 538 -6663 572
rect -6495 538 -6479 572
rect -6679 500 -6479 538
rect -6421 572 -6221 588
rect -6421 538 -6405 572
rect -6237 538 -6221 572
rect -6421 500 -6221 538
rect -6163 572 -5963 588
rect -6163 538 -6147 572
rect -5979 538 -5963 572
rect -6163 500 -5963 538
rect -5905 572 -5705 588
rect -5905 538 -5889 572
rect -5721 538 -5705 572
rect -5905 500 -5705 538
rect -5647 572 -5447 588
rect -5647 538 -5631 572
rect -5463 538 -5447 572
rect -5647 500 -5447 538
rect -5389 572 -5189 588
rect -5389 538 -5373 572
rect -5205 538 -5189 572
rect -5389 500 -5189 538
rect -5131 572 -4931 588
rect -5131 538 -5115 572
rect -4947 538 -4931 572
rect -5131 500 -4931 538
rect -4873 572 -4673 588
rect -4873 538 -4857 572
rect -4689 538 -4673 572
rect -4873 500 -4673 538
rect -4615 572 -4415 588
rect -4615 538 -4599 572
rect -4431 538 -4415 572
rect -4615 500 -4415 538
rect -4357 572 -4157 588
rect -4357 538 -4341 572
rect -4173 538 -4157 572
rect -4357 500 -4157 538
rect -4099 572 -3899 588
rect -4099 538 -4083 572
rect -3915 538 -3899 572
rect -4099 500 -3899 538
rect -3841 572 -3641 588
rect -3841 538 -3825 572
rect -3657 538 -3641 572
rect -3841 500 -3641 538
rect -3583 572 -3383 588
rect -3583 538 -3567 572
rect -3399 538 -3383 572
rect -3583 500 -3383 538
rect -3325 572 -3125 588
rect -3325 538 -3309 572
rect -3141 538 -3125 572
rect -3325 500 -3125 538
rect -3067 572 -2867 588
rect -3067 538 -3051 572
rect -2883 538 -2867 572
rect -3067 500 -2867 538
rect -2809 572 -2609 588
rect -2809 538 -2793 572
rect -2625 538 -2609 572
rect -2809 500 -2609 538
rect -2551 572 -2351 588
rect -2551 538 -2535 572
rect -2367 538 -2351 572
rect -2551 500 -2351 538
rect -2293 572 -2093 588
rect -2293 538 -2277 572
rect -2109 538 -2093 572
rect -2293 500 -2093 538
rect -2035 572 -1835 588
rect -2035 538 -2019 572
rect -1851 538 -1835 572
rect -2035 500 -1835 538
rect -1777 572 -1577 588
rect -1777 538 -1761 572
rect -1593 538 -1577 572
rect -1777 500 -1577 538
rect -1519 572 -1319 588
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1519 500 -1319 538
rect -1261 572 -1061 588
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1261 500 -1061 538
rect -1003 572 -803 588
rect -1003 538 -987 572
rect -819 538 -803 572
rect -1003 500 -803 538
rect -745 572 -545 588
rect -745 538 -729 572
rect -561 538 -545 572
rect -745 500 -545 538
rect -487 572 -287 588
rect -487 538 -471 572
rect -303 538 -287 572
rect -487 500 -287 538
rect -229 572 -29 588
rect -229 538 -213 572
rect -45 538 -29 572
rect -229 500 -29 538
rect 29 572 229 588
rect 29 538 45 572
rect 213 538 229 572
rect 29 500 229 538
rect 287 572 487 588
rect 287 538 303 572
rect 471 538 487 572
rect 287 500 487 538
rect 545 572 745 588
rect 545 538 561 572
rect 729 538 745 572
rect 545 500 745 538
rect 803 572 1003 588
rect 803 538 819 572
rect 987 538 1003 572
rect 803 500 1003 538
rect 1061 572 1261 588
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1061 500 1261 538
rect 1319 572 1519 588
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1319 500 1519 538
rect 1577 572 1777 588
rect 1577 538 1593 572
rect 1761 538 1777 572
rect 1577 500 1777 538
rect 1835 572 2035 588
rect 1835 538 1851 572
rect 2019 538 2035 572
rect 1835 500 2035 538
rect 2093 572 2293 588
rect 2093 538 2109 572
rect 2277 538 2293 572
rect 2093 500 2293 538
rect 2351 572 2551 588
rect 2351 538 2367 572
rect 2535 538 2551 572
rect 2351 500 2551 538
rect 2609 572 2809 588
rect 2609 538 2625 572
rect 2793 538 2809 572
rect 2609 500 2809 538
rect 2867 572 3067 588
rect 2867 538 2883 572
rect 3051 538 3067 572
rect 2867 500 3067 538
rect 3125 572 3325 588
rect 3125 538 3141 572
rect 3309 538 3325 572
rect 3125 500 3325 538
rect 3383 572 3583 588
rect 3383 538 3399 572
rect 3567 538 3583 572
rect 3383 500 3583 538
rect 3641 572 3841 588
rect 3641 538 3657 572
rect 3825 538 3841 572
rect 3641 500 3841 538
rect 3899 572 4099 588
rect 3899 538 3915 572
rect 4083 538 4099 572
rect 3899 500 4099 538
rect 4157 572 4357 588
rect 4157 538 4173 572
rect 4341 538 4357 572
rect 4157 500 4357 538
rect 4415 572 4615 588
rect 4415 538 4431 572
rect 4599 538 4615 572
rect 4415 500 4615 538
rect 4673 572 4873 588
rect 4673 538 4689 572
rect 4857 538 4873 572
rect 4673 500 4873 538
rect 4931 572 5131 588
rect 4931 538 4947 572
rect 5115 538 5131 572
rect 4931 500 5131 538
rect 5189 572 5389 588
rect 5189 538 5205 572
rect 5373 538 5389 572
rect 5189 500 5389 538
rect 5447 572 5647 588
rect 5447 538 5463 572
rect 5631 538 5647 572
rect 5447 500 5647 538
rect 5705 572 5905 588
rect 5705 538 5721 572
rect 5889 538 5905 572
rect 5705 500 5905 538
rect 5963 572 6163 588
rect 5963 538 5979 572
rect 6147 538 6163 572
rect 5963 500 6163 538
rect 6221 572 6421 588
rect 6221 538 6237 572
rect 6405 538 6421 572
rect 6221 500 6421 538
rect 6479 572 6679 588
rect 6479 538 6495 572
rect 6663 538 6679 572
rect 6479 500 6679 538
rect -6679 -538 -6479 -500
rect -6679 -572 -6663 -538
rect -6495 -572 -6479 -538
rect -6679 -588 -6479 -572
rect -6421 -538 -6221 -500
rect -6421 -572 -6405 -538
rect -6237 -572 -6221 -538
rect -6421 -588 -6221 -572
rect -6163 -538 -5963 -500
rect -6163 -572 -6147 -538
rect -5979 -572 -5963 -538
rect -6163 -588 -5963 -572
rect -5905 -538 -5705 -500
rect -5905 -572 -5889 -538
rect -5721 -572 -5705 -538
rect -5905 -588 -5705 -572
rect -5647 -538 -5447 -500
rect -5647 -572 -5631 -538
rect -5463 -572 -5447 -538
rect -5647 -588 -5447 -572
rect -5389 -538 -5189 -500
rect -5389 -572 -5373 -538
rect -5205 -572 -5189 -538
rect -5389 -588 -5189 -572
rect -5131 -538 -4931 -500
rect -5131 -572 -5115 -538
rect -4947 -572 -4931 -538
rect -5131 -588 -4931 -572
rect -4873 -538 -4673 -500
rect -4873 -572 -4857 -538
rect -4689 -572 -4673 -538
rect -4873 -588 -4673 -572
rect -4615 -538 -4415 -500
rect -4615 -572 -4599 -538
rect -4431 -572 -4415 -538
rect -4615 -588 -4415 -572
rect -4357 -538 -4157 -500
rect -4357 -572 -4341 -538
rect -4173 -572 -4157 -538
rect -4357 -588 -4157 -572
rect -4099 -538 -3899 -500
rect -4099 -572 -4083 -538
rect -3915 -572 -3899 -538
rect -4099 -588 -3899 -572
rect -3841 -538 -3641 -500
rect -3841 -572 -3825 -538
rect -3657 -572 -3641 -538
rect -3841 -588 -3641 -572
rect -3583 -538 -3383 -500
rect -3583 -572 -3567 -538
rect -3399 -572 -3383 -538
rect -3583 -588 -3383 -572
rect -3325 -538 -3125 -500
rect -3325 -572 -3309 -538
rect -3141 -572 -3125 -538
rect -3325 -588 -3125 -572
rect -3067 -538 -2867 -500
rect -3067 -572 -3051 -538
rect -2883 -572 -2867 -538
rect -3067 -588 -2867 -572
rect -2809 -538 -2609 -500
rect -2809 -572 -2793 -538
rect -2625 -572 -2609 -538
rect -2809 -588 -2609 -572
rect -2551 -538 -2351 -500
rect -2551 -572 -2535 -538
rect -2367 -572 -2351 -538
rect -2551 -588 -2351 -572
rect -2293 -538 -2093 -500
rect -2293 -572 -2277 -538
rect -2109 -572 -2093 -538
rect -2293 -588 -2093 -572
rect -2035 -538 -1835 -500
rect -2035 -572 -2019 -538
rect -1851 -572 -1835 -538
rect -2035 -588 -1835 -572
rect -1777 -538 -1577 -500
rect -1777 -572 -1761 -538
rect -1593 -572 -1577 -538
rect -1777 -588 -1577 -572
rect -1519 -538 -1319 -500
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1519 -588 -1319 -572
rect -1261 -538 -1061 -500
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1261 -588 -1061 -572
rect -1003 -538 -803 -500
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -1003 -588 -803 -572
rect -745 -538 -545 -500
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -745 -588 -545 -572
rect -487 -538 -287 -500
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -487 -588 -287 -572
rect -229 -538 -29 -500
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect -229 -588 -29 -572
rect 29 -538 229 -500
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 29 -588 229 -572
rect 287 -538 487 -500
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 287 -588 487 -572
rect 545 -538 745 -500
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 545 -588 745 -572
rect 803 -538 1003 -500
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 803 -588 1003 -572
rect 1061 -538 1261 -500
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1061 -588 1261 -572
rect 1319 -538 1519 -500
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1319 -588 1519 -572
rect 1577 -538 1777 -500
rect 1577 -572 1593 -538
rect 1761 -572 1777 -538
rect 1577 -588 1777 -572
rect 1835 -538 2035 -500
rect 1835 -572 1851 -538
rect 2019 -572 2035 -538
rect 1835 -588 2035 -572
rect 2093 -538 2293 -500
rect 2093 -572 2109 -538
rect 2277 -572 2293 -538
rect 2093 -588 2293 -572
rect 2351 -538 2551 -500
rect 2351 -572 2367 -538
rect 2535 -572 2551 -538
rect 2351 -588 2551 -572
rect 2609 -538 2809 -500
rect 2609 -572 2625 -538
rect 2793 -572 2809 -538
rect 2609 -588 2809 -572
rect 2867 -538 3067 -500
rect 2867 -572 2883 -538
rect 3051 -572 3067 -538
rect 2867 -588 3067 -572
rect 3125 -538 3325 -500
rect 3125 -572 3141 -538
rect 3309 -572 3325 -538
rect 3125 -588 3325 -572
rect 3383 -538 3583 -500
rect 3383 -572 3399 -538
rect 3567 -572 3583 -538
rect 3383 -588 3583 -572
rect 3641 -538 3841 -500
rect 3641 -572 3657 -538
rect 3825 -572 3841 -538
rect 3641 -588 3841 -572
rect 3899 -538 4099 -500
rect 3899 -572 3915 -538
rect 4083 -572 4099 -538
rect 3899 -588 4099 -572
rect 4157 -538 4357 -500
rect 4157 -572 4173 -538
rect 4341 -572 4357 -538
rect 4157 -588 4357 -572
rect 4415 -538 4615 -500
rect 4415 -572 4431 -538
rect 4599 -572 4615 -538
rect 4415 -588 4615 -572
rect 4673 -538 4873 -500
rect 4673 -572 4689 -538
rect 4857 -572 4873 -538
rect 4673 -588 4873 -572
rect 4931 -538 5131 -500
rect 4931 -572 4947 -538
rect 5115 -572 5131 -538
rect 4931 -588 5131 -572
rect 5189 -538 5389 -500
rect 5189 -572 5205 -538
rect 5373 -572 5389 -538
rect 5189 -588 5389 -572
rect 5447 -538 5647 -500
rect 5447 -572 5463 -538
rect 5631 -572 5647 -538
rect 5447 -588 5647 -572
rect 5705 -538 5905 -500
rect 5705 -572 5721 -538
rect 5889 -572 5905 -538
rect 5705 -588 5905 -572
rect 5963 -538 6163 -500
rect 5963 -572 5979 -538
rect 6147 -572 6163 -538
rect 5963 -588 6163 -572
rect 6221 -538 6421 -500
rect 6221 -572 6237 -538
rect 6405 -572 6421 -538
rect 6221 -588 6421 -572
rect 6479 -538 6679 -500
rect 6479 -572 6495 -538
rect 6663 -572 6679 -538
rect 6479 -588 6679 -572
<< polycont >>
rect -6663 538 -6495 572
rect -6405 538 -6237 572
rect -6147 538 -5979 572
rect -5889 538 -5721 572
rect -5631 538 -5463 572
rect -5373 538 -5205 572
rect -5115 538 -4947 572
rect -4857 538 -4689 572
rect -4599 538 -4431 572
rect -4341 538 -4173 572
rect -4083 538 -3915 572
rect -3825 538 -3657 572
rect -3567 538 -3399 572
rect -3309 538 -3141 572
rect -3051 538 -2883 572
rect -2793 538 -2625 572
rect -2535 538 -2367 572
rect -2277 538 -2109 572
rect -2019 538 -1851 572
rect -1761 538 -1593 572
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect 1593 538 1761 572
rect 1851 538 2019 572
rect 2109 538 2277 572
rect 2367 538 2535 572
rect 2625 538 2793 572
rect 2883 538 3051 572
rect 3141 538 3309 572
rect 3399 538 3567 572
rect 3657 538 3825 572
rect 3915 538 4083 572
rect 4173 538 4341 572
rect 4431 538 4599 572
rect 4689 538 4857 572
rect 4947 538 5115 572
rect 5205 538 5373 572
rect 5463 538 5631 572
rect 5721 538 5889 572
rect 5979 538 6147 572
rect 6237 538 6405 572
rect 6495 538 6663 572
rect -6663 -572 -6495 -538
rect -6405 -572 -6237 -538
rect -6147 -572 -5979 -538
rect -5889 -572 -5721 -538
rect -5631 -572 -5463 -538
rect -5373 -572 -5205 -538
rect -5115 -572 -4947 -538
rect -4857 -572 -4689 -538
rect -4599 -572 -4431 -538
rect -4341 -572 -4173 -538
rect -4083 -572 -3915 -538
rect -3825 -572 -3657 -538
rect -3567 -572 -3399 -538
rect -3309 -572 -3141 -538
rect -3051 -572 -2883 -538
rect -2793 -572 -2625 -538
rect -2535 -572 -2367 -538
rect -2277 -572 -2109 -538
rect -2019 -572 -1851 -538
rect -1761 -572 -1593 -538
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
rect 1593 -572 1761 -538
rect 1851 -572 2019 -538
rect 2109 -572 2277 -538
rect 2367 -572 2535 -538
rect 2625 -572 2793 -538
rect 2883 -572 3051 -538
rect 3141 -572 3309 -538
rect 3399 -572 3567 -538
rect 3657 -572 3825 -538
rect 3915 -572 4083 -538
rect 4173 -572 4341 -538
rect 4431 -572 4599 -538
rect 4689 -572 4857 -538
rect 4947 -572 5115 -538
rect 5205 -572 5373 -538
rect 5463 -572 5631 -538
rect 5721 -572 5889 -538
rect 5979 -572 6147 -538
rect 6237 -572 6405 -538
rect 6495 -572 6663 -538
<< locali >>
rect -6861 676 -6765 710
rect 6765 676 6861 710
rect -6861 614 -6827 676
rect 6827 614 6861 676
rect -6679 538 -6663 572
rect -6495 538 -6479 572
rect -6421 538 -6405 572
rect -6237 538 -6221 572
rect -6163 538 -6147 572
rect -5979 538 -5963 572
rect -5905 538 -5889 572
rect -5721 538 -5705 572
rect -5647 538 -5631 572
rect -5463 538 -5447 572
rect -5389 538 -5373 572
rect -5205 538 -5189 572
rect -5131 538 -5115 572
rect -4947 538 -4931 572
rect -4873 538 -4857 572
rect -4689 538 -4673 572
rect -4615 538 -4599 572
rect -4431 538 -4415 572
rect -4357 538 -4341 572
rect -4173 538 -4157 572
rect -4099 538 -4083 572
rect -3915 538 -3899 572
rect -3841 538 -3825 572
rect -3657 538 -3641 572
rect -3583 538 -3567 572
rect -3399 538 -3383 572
rect -3325 538 -3309 572
rect -3141 538 -3125 572
rect -3067 538 -3051 572
rect -2883 538 -2867 572
rect -2809 538 -2793 572
rect -2625 538 -2609 572
rect -2551 538 -2535 572
rect -2367 538 -2351 572
rect -2293 538 -2277 572
rect -2109 538 -2093 572
rect -2035 538 -2019 572
rect -1851 538 -1835 572
rect -1777 538 -1761 572
rect -1593 538 -1577 572
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1003 538 -987 572
rect -819 538 -803 572
rect -745 538 -729 572
rect -561 538 -545 572
rect -487 538 -471 572
rect -303 538 -287 572
rect -229 538 -213 572
rect -45 538 -29 572
rect 29 538 45 572
rect 213 538 229 572
rect 287 538 303 572
rect 471 538 487 572
rect 545 538 561 572
rect 729 538 745 572
rect 803 538 819 572
rect 987 538 1003 572
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1577 538 1593 572
rect 1761 538 1777 572
rect 1835 538 1851 572
rect 2019 538 2035 572
rect 2093 538 2109 572
rect 2277 538 2293 572
rect 2351 538 2367 572
rect 2535 538 2551 572
rect 2609 538 2625 572
rect 2793 538 2809 572
rect 2867 538 2883 572
rect 3051 538 3067 572
rect 3125 538 3141 572
rect 3309 538 3325 572
rect 3383 538 3399 572
rect 3567 538 3583 572
rect 3641 538 3657 572
rect 3825 538 3841 572
rect 3899 538 3915 572
rect 4083 538 4099 572
rect 4157 538 4173 572
rect 4341 538 4357 572
rect 4415 538 4431 572
rect 4599 538 4615 572
rect 4673 538 4689 572
rect 4857 538 4873 572
rect 4931 538 4947 572
rect 5115 538 5131 572
rect 5189 538 5205 572
rect 5373 538 5389 572
rect 5447 538 5463 572
rect 5631 538 5647 572
rect 5705 538 5721 572
rect 5889 538 5905 572
rect 5963 538 5979 572
rect 6147 538 6163 572
rect 6221 538 6237 572
rect 6405 538 6421 572
rect 6479 538 6495 572
rect 6663 538 6679 572
rect -6725 488 -6691 504
rect -6725 -504 -6691 -488
rect -6467 488 -6433 504
rect -6467 -504 -6433 -488
rect -6209 488 -6175 504
rect -6209 -504 -6175 -488
rect -5951 488 -5917 504
rect -5951 -504 -5917 -488
rect -5693 488 -5659 504
rect -5693 -504 -5659 -488
rect -5435 488 -5401 504
rect -5435 -504 -5401 -488
rect -5177 488 -5143 504
rect -5177 -504 -5143 -488
rect -4919 488 -4885 504
rect -4919 -504 -4885 -488
rect -4661 488 -4627 504
rect -4661 -504 -4627 -488
rect -4403 488 -4369 504
rect -4403 -504 -4369 -488
rect -4145 488 -4111 504
rect -4145 -504 -4111 -488
rect -3887 488 -3853 504
rect -3887 -504 -3853 -488
rect -3629 488 -3595 504
rect -3629 -504 -3595 -488
rect -3371 488 -3337 504
rect -3371 -504 -3337 -488
rect -3113 488 -3079 504
rect -3113 -504 -3079 -488
rect -2855 488 -2821 504
rect -2855 -504 -2821 -488
rect -2597 488 -2563 504
rect -2597 -504 -2563 -488
rect -2339 488 -2305 504
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect 2305 488 2339 504
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -504 2597 -488
rect 2821 488 2855 504
rect 2821 -504 2855 -488
rect 3079 488 3113 504
rect 3079 -504 3113 -488
rect 3337 488 3371 504
rect 3337 -504 3371 -488
rect 3595 488 3629 504
rect 3595 -504 3629 -488
rect 3853 488 3887 504
rect 3853 -504 3887 -488
rect 4111 488 4145 504
rect 4111 -504 4145 -488
rect 4369 488 4403 504
rect 4369 -504 4403 -488
rect 4627 488 4661 504
rect 4627 -504 4661 -488
rect 4885 488 4919 504
rect 4885 -504 4919 -488
rect 5143 488 5177 504
rect 5143 -504 5177 -488
rect 5401 488 5435 504
rect 5401 -504 5435 -488
rect 5659 488 5693 504
rect 5659 -504 5693 -488
rect 5917 488 5951 504
rect 5917 -504 5951 -488
rect 6175 488 6209 504
rect 6175 -504 6209 -488
rect 6433 488 6467 504
rect 6433 -504 6467 -488
rect 6691 488 6725 504
rect 6691 -504 6725 -488
rect -6679 -572 -6663 -538
rect -6495 -572 -6479 -538
rect -6421 -572 -6405 -538
rect -6237 -572 -6221 -538
rect -6163 -572 -6147 -538
rect -5979 -572 -5963 -538
rect -5905 -572 -5889 -538
rect -5721 -572 -5705 -538
rect -5647 -572 -5631 -538
rect -5463 -572 -5447 -538
rect -5389 -572 -5373 -538
rect -5205 -572 -5189 -538
rect -5131 -572 -5115 -538
rect -4947 -572 -4931 -538
rect -4873 -572 -4857 -538
rect -4689 -572 -4673 -538
rect -4615 -572 -4599 -538
rect -4431 -572 -4415 -538
rect -4357 -572 -4341 -538
rect -4173 -572 -4157 -538
rect -4099 -572 -4083 -538
rect -3915 -572 -3899 -538
rect -3841 -572 -3825 -538
rect -3657 -572 -3641 -538
rect -3583 -572 -3567 -538
rect -3399 -572 -3383 -538
rect -3325 -572 -3309 -538
rect -3141 -572 -3125 -538
rect -3067 -572 -3051 -538
rect -2883 -572 -2867 -538
rect -2809 -572 -2793 -538
rect -2625 -572 -2609 -538
rect -2551 -572 -2535 -538
rect -2367 -572 -2351 -538
rect -2293 -572 -2277 -538
rect -2109 -572 -2093 -538
rect -2035 -572 -2019 -538
rect -1851 -572 -1835 -538
rect -1777 -572 -1761 -538
rect -1593 -572 -1577 -538
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1577 -572 1593 -538
rect 1761 -572 1777 -538
rect 1835 -572 1851 -538
rect 2019 -572 2035 -538
rect 2093 -572 2109 -538
rect 2277 -572 2293 -538
rect 2351 -572 2367 -538
rect 2535 -572 2551 -538
rect 2609 -572 2625 -538
rect 2793 -572 2809 -538
rect 2867 -572 2883 -538
rect 3051 -572 3067 -538
rect 3125 -572 3141 -538
rect 3309 -572 3325 -538
rect 3383 -572 3399 -538
rect 3567 -572 3583 -538
rect 3641 -572 3657 -538
rect 3825 -572 3841 -538
rect 3899 -572 3915 -538
rect 4083 -572 4099 -538
rect 4157 -572 4173 -538
rect 4341 -572 4357 -538
rect 4415 -572 4431 -538
rect 4599 -572 4615 -538
rect 4673 -572 4689 -538
rect 4857 -572 4873 -538
rect 4931 -572 4947 -538
rect 5115 -572 5131 -538
rect 5189 -572 5205 -538
rect 5373 -572 5389 -538
rect 5447 -572 5463 -538
rect 5631 -572 5647 -538
rect 5705 -572 5721 -538
rect 5889 -572 5905 -538
rect 5963 -572 5979 -538
rect 6147 -572 6163 -538
rect 6221 -572 6237 -538
rect 6405 -572 6421 -538
rect 6479 -572 6495 -538
rect 6663 -572 6679 -538
rect -6861 -676 -6827 -614
rect 6827 -676 6861 -614
rect -6861 -710 -6765 -676
rect 6765 -710 6861 -676
<< viali >>
rect -6663 538 -6495 572
rect -6405 538 -6237 572
rect -6147 538 -5979 572
rect -5889 538 -5721 572
rect -5631 538 -5463 572
rect -5373 538 -5205 572
rect -5115 538 -4947 572
rect -4857 538 -4689 572
rect -4599 538 -4431 572
rect -4341 538 -4173 572
rect -4083 538 -3915 572
rect -3825 538 -3657 572
rect -3567 538 -3399 572
rect -3309 538 -3141 572
rect -3051 538 -2883 572
rect -2793 538 -2625 572
rect -2535 538 -2367 572
rect -2277 538 -2109 572
rect -2019 538 -1851 572
rect -1761 538 -1593 572
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect 1593 538 1761 572
rect 1851 538 2019 572
rect 2109 538 2277 572
rect 2367 538 2535 572
rect 2625 538 2793 572
rect 2883 538 3051 572
rect 3141 538 3309 572
rect 3399 538 3567 572
rect 3657 538 3825 572
rect 3915 538 4083 572
rect 4173 538 4341 572
rect 4431 538 4599 572
rect 4689 538 4857 572
rect 4947 538 5115 572
rect 5205 538 5373 572
rect 5463 538 5631 572
rect 5721 538 5889 572
rect 5979 538 6147 572
rect 6237 538 6405 572
rect 6495 538 6663 572
rect -6725 -488 -6691 488
rect -6467 -488 -6433 488
rect -6209 -488 -6175 488
rect -5951 -488 -5917 488
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect 5917 -488 5951 488
rect 6175 -488 6209 488
rect 6433 -488 6467 488
rect 6691 -488 6725 488
rect -6663 -572 -6495 -538
rect -6405 -572 -6237 -538
rect -6147 -572 -5979 -538
rect -5889 -572 -5721 -538
rect -5631 -572 -5463 -538
rect -5373 -572 -5205 -538
rect -5115 -572 -4947 -538
rect -4857 -572 -4689 -538
rect -4599 -572 -4431 -538
rect -4341 -572 -4173 -538
rect -4083 -572 -3915 -538
rect -3825 -572 -3657 -538
rect -3567 -572 -3399 -538
rect -3309 -572 -3141 -538
rect -3051 -572 -2883 -538
rect -2793 -572 -2625 -538
rect -2535 -572 -2367 -538
rect -2277 -572 -2109 -538
rect -2019 -572 -1851 -538
rect -1761 -572 -1593 -538
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
rect 1593 -572 1761 -538
rect 1851 -572 2019 -538
rect 2109 -572 2277 -538
rect 2367 -572 2535 -538
rect 2625 -572 2793 -538
rect 2883 -572 3051 -538
rect 3141 -572 3309 -538
rect 3399 -572 3567 -538
rect 3657 -572 3825 -538
rect 3915 -572 4083 -538
rect 4173 -572 4341 -538
rect 4431 -572 4599 -538
rect 4689 -572 4857 -538
rect 4947 -572 5115 -538
rect 5205 -572 5373 -538
rect 5463 -572 5631 -538
rect 5721 -572 5889 -538
rect 5979 -572 6147 -538
rect 6237 -572 6405 -538
rect 6495 -572 6663 -538
<< metal1 >>
rect -6675 572 -6483 578
rect -6675 538 -6663 572
rect -6495 538 -6483 572
rect -6675 532 -6483 538
rect -6417 572 -6225 578
rect -6417 538 -6405 572
rect -6237 538 -6225 572
rect -6417 532 -6225 538
rect -6159 572 -5967 578
rect -6159 538 -6147 572
rect -5979 538 -5967 572
rect -6159 532 -5967 538
rect -5901 572 -5709 578
rect -5901 538 -5889 572
rect -5721 538 -5709 572
rect -5901 532 -5709 538
rect -5643 572 -5451 578
rect -5643 538 -5631 572
rect -5463 538 -5451 572
rect -5643 532 -5451 538
rect -5385 572 -5193 578
rect -5385 538 -5373 572
rect -5205 538 -5193 572
rect -5385 532 -5193 538
rect -5127 572 -4935 578
rect -5127 538 -5115 572
rect -4947 538 -4935 572
rect -5127 532 -4935 538
rect -4869 572 -4677 578
rect -4869 538 -4857 572
rect -4689 538 -4677 572
rect -4869 532 -4677 538
rect -4611 572 -4419 578
rect -4611 538 -4599 572
rect -4431 538 -4419 572
rect -4611 532 -4419 538
rect -4353 572 -4161 578
rect -4353 538 -4341 572
rect -4173 538 -4161 572
rect -4353 532 -4161 538
rect -4095 572 -3903 578
rect -4095 538 -4083 572
rect -3915 538 -3903 572
rect -4095 532 -3903 538
rect -3837 572 -3645 578
rect -3837 538 -3825 572
rect -3657 538 -3645 572
rect -3837 532 -3645 538
rect -3579 572 -3387 578
rect -3579 538 -3567 572
rect -3399 538 -3387 572
rect -3579 532 -3387 538
rect -3321 572 -3129 578
rect -3321 538 -3309 572
rect -3141 538 -3129 572
rect -3321 532 -3129 538
rect -3063 572 -2871 578
rect -3063 538 -3051 572
rect -2883 538 -2871 572
rect -3063 532 -2871 538
rect -2805 572 -2613 578
rect -2805 538 -2793 572
rect -2625 538 -2613 572
rect -2805 532 -2613 538
rect -2547 572 -2355 578
rect -2547 538 -2535 572
rect -2367 538 -2355 572
rect -2547 532 -2355 538
rect -2289 572 -2097 578
rect -2289 538 -2277 572
rect -2109 538 -2097 572
rect -2289 532 -2097 538
rect -2031 572 -1839 578
rect -2031 538 -2019 572
rect -1851 538 -1839 572
rect -2031 532 -1839 538
rect -1773 572 -1581 578
rect -1773 538 -1761 572
rect -1593 538 -1581 572
rect -1773 532 -1581 538
rect -1515 572 -1323 578
rect -1515 538 -1503 572
rect -1335 538 -1323 572
rect -1515 532 -1323 538
rect -1257 572 -1065 578
rect -1257 538 -1245 572
rect -1077 538 -1065 572
rect -1257 532 -1065 538
rect -999 572 -807 578
rect -999 538 -987 572
rect -819 538 -807 572
rect -999 532 -807 538
rect -741 572 -549 578
rect -741 538 -729 572
rect -561 538 -549 572
rect -741 532 -549 538
rect -483 572 -291 578
rect -483 538 -471 572
rect -303 538 -291 572
rect -483 532 -291 538
rect -225 572 -33 578
rect -225 538 -213 572
rect -45 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 45 572
rect 213 538 225 572
rect 33 532 225 538
rect 291 572 483 578
rect 291 538 303 572
rect 471 538 483 572
rect 291 532 483 538
rect 549 572 741 578
rect 549 538 561 572
rect 729 538 741 572
rect 549 532 741 538
rect 807 572 999 578
rect 807 538 819 572
rect 987 538 999 572
rect 807 532 999 538
rect 1065 572 1257 578
rect 1065 538 1077 572
rect 1245 538 1257 572
rect 1065 532 1257 538
rect 1323 572 1515 578
rect 1323 538 1335 572
rect 1503 538 1515 572
rect 1323 532 1515 538
rect 1581 572 1773 578
rect 1581 538 1593 572
rect 1761 538 1773 572
rect 1581 532 1773 538
rect 1839 572 2031 578
rect 1839 538 1851 572
rect 2019 538 2031 572
rect 1839 532 2031 538
rect 2097 572 2289 578
rect 2097 538 2109 572
rect 2277 538 2289 572
rect 2097 532 2289 538
rect 2355 572 2547 578
rect 2355 538 2367 572
rect 2535 538 2547 572
rect 2355 532 2547 538
rect 2613 572 2805 578
rect 2613 538 2625 572
rect 2793 538 2805 572
rect 2613 532 2805 538
rect 2871 572 3063 578
rect 2871 538 2883 572
rect 3051 538 3063 572
rect 2871 532 3063 538
rect 3129 572 3321 578
rect 3129 538 3141 572
rect 3309 538 3321 572
rect 3129 532 3321 538
rect 3387 572 3579 578
rect 3387 538 3399 572
rect 3567 538 3579 572
rect 3387 532 3579 538
rect 3645 572 3837 578
rect 3645 538 3657 572
rect 3825 538 3837 572
rect 3645 532 3837 538
rect 3903 572 4095 578
rect 3903 538 3915 572
rect 4083 538 4095 572
rect 3903 532 4095 538
rect 4161 572 4353 578
rect 4161 538 4173 572
rect 4341 538 4353 572
rect 4161 532 4353 538
rect 4419 572 4611 578
rect 4419 538 4431 572
rect 4599 538 4611 572
rect 4419 532 4611 538
rect 4677 572 4869 578
rect 4677 538 4689 572
rect 4857 538 4869 572
rect 4677 532 4869 538
rect 4935 572 5127 578
rect 4935 538 4947 572
rect 5115 538 5127 572
rect 4935 532 5127 538
rect 5193 572 5385 578
rect 5193 538 5205 572
rect 5373 538 5385 572
rect 5193 532 5385 538
rect 5451 572 5643 578
rect 5451 538 5463 572
rect 5631 538 5643 572
rect 5451 532 5643 538
rect 5709 572 5901 578
rect 5709 538 5721 572
rect 5889 538 5901 572
rect 5709 532 5901 538
rect 5967 572 6159 578
rect 5967 538 5979 572
rect 6147 538 6159 572
rect 5967 532 6159 538
rect 6225 572 6417 578
rect 6225 538 6237 572
rect 6405 538 6417 572
rect 6225 532 6417 538
rect 6483 572 6675 578
rect 6483 538 6495 572
rect 6663 538 6675 572
rect 6483 532 6675 538
rect -6731 488 -6685 500
rect -6731 -488 -6725 488
rect -6691 -488 -6685 488
rect -6731 -500 -6685 -488
rect -6473 488 -6427 500
rect -6473 -488 -6467 488
rect -6433 -488 -6427 488
rect -6473 -500 -6427 -488
rect -6215 488 -6169 500
rect -6215 -488 -6209 488
rect -6175 -488 -6169 488
rect -6215 -500 -6169 -488
rect -5957 488 -5911 500
rect -5957 -488 -5951 488
rect -5917 -488 -5911 488
rect -5957 -500 -5911 -488
rect -5699 488 -5653 500
rect -5699 -488 -5693 488
rect -5659 -488 -5653 488
rect -5699 -500 -5653 -488
rect -5441 488 -5395 500
rect -5441 -488 -5435 488
rect -5401 -488 -5395 488
rect -5441 -500 -5395 -488
rect -5183 488 -5137 500
rect -5183 -488 -5177 488
rect -5143 -488 -5137 488
rect -5183 -500 -5137 -488
rect -4925 488 -4879 500
rect -4925 -488 -4919 488
rect -4885 -488 -4879 488
rect -4925 -500 -4879 -488
rect -4667 488 -4621 500
rect -4667 -488 -4661 488
rect -4627 -488 -4621 488
rect -4667 -500 -4621 -488
rect -4409 488 -4363 500
rect -4409 -488 -4403 488
rect -4369 -488 -4363 488
rect -4409 -500 -4363 -488
rect -4151 488 -4105 500
rect -4151 -488 -4145 488
rect -4111 -488 -4105 488
rect -4151 -500 -4105 -488
rect -3893 488 -3847 500
rect -3893 -488 -3887 488
rect -3853 -488 -3847 488
rect -3893 -500 -3847 -488
rect -3635 488 -3589 500
rect -3635 -488 -3629 488
rect -3595 -488 -3589 488
rect -3635 -500 -3589 -488
rect -3377 488 -3331 500
rect -3377 -488 -3371 488
rect -3337 -488 -3331 488
rect -3377 -500 -3331 -488
rect -3119 488 -3073 500
rect -3119 -488 -3113 488
rect -3079 -488 -3073 488
rect -3119 -500 -3073 -488
rect -2861 488 -2815 500
rect -2861 -488 -2855 488
rect -2821 -488 -2815 488
rect -2861 -500 -2815 -488
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect 2815 488 2861 500
rect 2815 -488 2821 488
rect 2855 -488 2861 488
rect 2815 -500 2861 -488
rect 3073 488 3119 500
rect 3073 -488 3079 488
rect 3113 -488 3119 488
rect 3073 -500 3119 -488
rect 3331 488 3377 500
rect 3331 -488 3337 488
rect 3371 -488 3377 488
rect 3331 -500 3377 -488
rect 3589 488 3635 500
rect 3589 -488 3595 488
rect 3629 -488 3635 488
rect 3589 -500 3635 -488
rect 3847 488 3893 500
rect 3847 -488 3853 488
rect 3887 -488 3893 488
rect 3847 -500 3893 -488
rect 4105 488 4151 500
rect 4105 -488 4111 488
rect 4145 -488 4151 488
rect 4105 -500 4151 -488
rect 4363 488 4409 500
rect 4363 -488 4369 488
rect 4403 -488 4409 488
rect 4363 -500 4409 -488
rect 4621 488 4667 500
rect 4621 -488 4627 488
rect 4661 -488 4667 488
rect 4621 -500 4667 -488
rect 4879 488 4925 500
rect 4879 -488 4885 488
rect 4919 -488 4925 488
rect 4879 -500 4925 -488
rect 5137 488 5183 500
rect 5137 -488 5143 488
rect 5177 -488 5183 488
rect 5137 -500 5183 -488
rect 5395 488 5441 500
rect 5395 -488 5401 488
rect 5435 -488 5441 488
rect 5395 -500 5441 -488
rect 5653 488 5699 500
rect 5653 -488 5659 488
rect 5693 -488 5699 488
rect 5653 -500 5699 -488
rect 5911 488 5957 500
rect 5911 -488 5917 488
rect 5951 -488 5957 488
rect 5911 -500 5957 -488
rect 6169 488 6215 500
rect 6169 -488 6175 488
rect 6209 -488 6215 488
rect 6169 -500 6215 -488
rect 6427 488 6473 500
rect 6427 -488 6433 488
rect 6467 -488 6473 488
rect 6427 -500 6473 -488
rect 6685 488 6731 500
rect 6685 -488 6691 488
rect 6725 -488 6731 488
rect 6685 -500 6731 -488
rect -6675 -538 -6483 -532
rect -6675 -572 -6663 -538
rect -6495 -572 -6483 -538
rect -6675 -578 -6483 -572
rect -6417 -538 -6225 -532
rect -6417 -572 -6405 -538
rect -6237 -572 -6225 -538
rect -6417 -578 -6225 -572
rect -6159 -538 -5967 -532
rect -6159 -572 -6147 -538
rect -5979 -572 -5967 -538
rect -6159 -578 -5967 -572
rect -5901 -538 -5709 -532
rect -5901 -572 -5889 -538
rect -5721 -572 -5709 -538
rect -5901 -578 -5709 -572
rect -5643 -538 -5451 -532
rect -5643 -572 -5631 -538
rect -5463 -572 -5451 -538
rect -5643 -578 -5451 -572
rect -5385 -538 -5193 -532
rect -5385 -572 -5373 -538
rect -5205 -572 -5193 -538
rect -5385 -578 -5193 -572
rect -5127 -538 -4935 -532
rect -5127 -572 -5115 -538
rect -4947 -572 -4935 -538
rect -5127 -578 -4935 -572
rect -4869 -538 -4677 -532
rect -4869 -572 -4857 -538
rect -4689 -572 -4677 -538
rect -4869 -578 -4677 -572
rect -4611 -538 -4419 -532
rect -4611 -572 -4599 -538
rect -4431 -572 -4419 -538
rect -4611 -578 -4419 -572
rect -4353 -538 -4161 -532
rect -4353 -572 -4341 -538
rect -4173 -572 -4161 -538
rect -4353 -578 -4161 -572
rect -4095 -538 -3903 -532
rect -4095 -572 -4083 -538
rect -3915 -572 -3903 -538
rect -4095 -578 -3903 -572
rect -3837 -538 -3645 -532
rect -3837 -572 -3825 -538
rect -3657 -572 -3645 -538
rect -3837 -578 -3645 -572
rect -3579 -538 -3387 -532
rect -3579 -572 -3567 -538
rect -3399 -572 -3387 -538
rect -3579 -578 -3387 -572
rect -3321 -538 -3129 -532
rect -3321 -572 -3309 -538
rect -3141 -572 -3129 -538
rect -3321 -578 -3129 -572
rect -3063 -538 -2871 -532
rect -3063 -572 -3051 -538
rect -2883 -572 -2871 -538
rect -3063 -578 -2871 -572
rect -2805 -538 -2613 -532
rect -2805 -572 -2793 -538
rect -2625 -572 -2613 -538
rect -2805 -578 -2613 -572
rect -2547 -538 -2355 -532
rect -2547 -572 -2535 -538
rect -2367 -572 -2355 -538
rect -2547 -578 -2355 -572
rect -2289 -538 -2097 -532
rect -2289 -572 -2277 -538
rect -2109 -572 -2097 -538
rect -2289 -578 -2097 -572
rect -2031 -538 -1839 -532
rect -2031 -572 -2019 -538
rect -1851 -572 -1839 -538
rect -2031 -578 -1839 -572
rect -1773 -538 -1581 -532
rect -1773 -572 -1761 -538
rect -1593 -572 -1581 -538
rect -1773 -578 -1581 -572
rect -1515 -538 -1323 -532
rect -1515 -572 -1503 -538
rect -1335 -572 -1323 -538
rect -1515 -578 -1323 -572
rect -1257 -538 -1065 -532
rect -1257 -572 -1245 -538
rect -1077 -572 -1065 -538
rect -1257 -578 -1065 -572
rect -999 -538 -807 -532
rect -999 -572 -987 -538
rect -819 -572 -807 -538
rect -999 -578 -807 -572
rect -741 -538 -549 -532
rect -741 -572 -729 -538
rect -561 -572 -549 -538
rect -741 -578 -549 -572
rect -483 -538 -291 -532
rect -483 -572 -471 -538
rect -303 -572 -291 -538
rect -483 -578 -291 -572
rect -225 -538 -33 -532
rect -225 -572 -213 -538
rect -45 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 45 -538
rect 213 -572 225 -538
rect 33 -578 225 -572
rect 291 -538 483 -532
rect 291 -572 303 -538
rect 471 -572 483 -538
rect 291 -578 483 -572
rect 549 -538 741 -532
rect 549 -572 561 -538
rect 729 -572 741 -538
rect 549 -578 741 -572
rect 807 -538 999 -532
rect 807 -572 819 -538
rect 987 -572 999 -538
rect 807 -578 999 -572
rect 1065 -538 1257 -532
rect 1065 -572 1077 -538
rect 1245 -572 1257 -538
rect 1065 -578 1257 -572
rect 1323 -538 1515 -532
rect 1323 -572 1335 -538
rect 1503 -572 1515 -538
rect 1323 -578 1515 -572
rect 1581 -538 1773 -532
rect 1581 -572 1593 -538
rect 1761 -572 1773 -538
rect 1581 -578 1773 -572
rect 1839 -538 2031 -532
rect 1839 -572 1851 -538
rect 2019 -572 2031 -538
rect 1839 -578 2031 -572
rect 2097 -538 2289 -532
rect 2097 -572 2109 -538
rect 2277 -572 2289 -538
rect 2097 -578 2289 -572
rect 2355 -538 2547 -532
rect 2355 -572 2367 -538
rect 2535 -572 2547 -538
rect 2355 -578 2547 -572
rect 2613 -538 2805 -532
rect 2613 -572 2625 -538
rect 2793 -572 2805 -538
rect 2613 -578 2805 -572
rect 2871 -538 3063 -532
rect 2871 -572 2883 -538
rect 3051 -572 3063 -538
rect 2871 -578 3063 -572
rect 3129 -538 3321 -532
rect 3129 -572 3141 -538
rect 3309 -572 3321 -538
rect 3129 -578 3321 -572
rect 3387 -538 3579 -532
rect 3387 -572 3399 -538
rect 3567 -572 3579 -538
rect 3387 -578 3579 -572
rect 3645 -538 3837 -532
rect 3645 -572 3657 -538
rect 3825 -572 3837 -538
rect 3645 -578 3837 -572
rect 3903 -538 4095 -532
rect 3903 -572 3915 -538
rect 4083 -572 4095 -538
rect 3903 -578 4095 -572
rect 4161 -538 4353 -532
rect 4161 -572 4173 -538
rect 4341 -572 4353 -538
rect 4161 -578 4353 -572
rect 4419 -538 4611 -532
rect 4419 -572 4431 -538
rect 4599 -572 4611 -538
rect 4419 -578 4611 -572
rect 4677 -538 4869 -532
rect 4677 -572 4689 -538
rect 4857 -572 4869 -538
rect 4677 -578 4869 -572
rect 4935 -538 5127 -532
rect 4935 -572 4947 -538
rect 5115 -572 5127 -538
rect 4935 -578 5127 -572
rect 5193 -538 5385 -532
rect 5193 -572 5205 -538
rect 5373 -572 5385 -538
rect 5193 -578 5385 -572
rect 5451 -538 5643 -532
rect 5451 -572 5463 -538
rect 5631 -572 5643 -538
rect 5451 -578 5643 -572
rect 5709 -538 5901 -532
rect 5709 -572 5721 -538
rect 5889 -572 5901 -538
rect 5709 -578 5901 -572
rect 5967 -538 6159 -532
rect 5967 -572 5979 -538
rect 6147 -572 6159 -538
rect 5967 -578 6159 -572
rect 6225 -538 6417 -532
rect 6225 -572 6237 -538
rect 6405 -572 6417 -538
rect 6225 -578 6417 -572
rect 6483 -538 6675 -532
rect 6483 -572 6495 -538
rect 6663 -572 6675 -538
rect 6483 -578 6675 -572
<< labels >>
rlabel mvpsubdiffcont 0 -693 0 -693 0 B
port 1 nsew
rlabel mvndiffc -6708 0 -6708 0 0 D0
port 2 nsew
rlabel polycont -6579 555 -6579 555 0 G0
port 3 nsew
rlabel mvndiffc -6450 0 -6450 0 0 S1
port 4 nsew
rlabel polycont -6321 555 -6321 555 0 G1
port 5 nsew
rlabel mvndiffc -6192 0 -6192 0 0 D2
port 6 nsew
rlabel polycont -6063 555 -6063 555 0 G2
port 7 nsew
rlabel mvndiffc -5934 0 -5934 0 0 S3
port 8 nsew
rlabel polycont -5805 555 -5805 555 0 G3
port 9 nsew
rlabel mvndiffc -5676 0 -5676 0 0 D4
port 10 nsew
rlabel polycont -5547 555 -5547 555 0 G4
port 11 nsew
rlabel mvndiffc -5418 0 -5418 0 0 S5
port 12 nsew
rlabel polycont -5289 555 -5289 555 0 G5
port 13 nsew
rlabel mvndiffc -5160 0 -5160 0 0 D6
port 14 nsew
rlabel polycont -5031 555 -5031 555 0 G6
port 15 nsew
rlabel mvndiffc -4902 0 -4902 0 0 S7
port 16 nsew
rlabel polycont -4773 555 -4773 555 0 G7
port 17 nsew
rlabel mvndiffc -4644 0 -4644 0 0 D8
port 18 nsew
rlabel polycont -4515 555 -4515 555 0 G8
port 19 nsew
rlabel mvndiffc -4386 0 -4386 0 0 S9
port 20 nsew
rlabel polycont -4257 555 -4257 555 0 G9
port 21 nsew
rlabel mvndiffc -4128 0 -4128 0 0 D10
port 22 nsew
rlabel polycont -3999 555 -3999 555 0 G10
port 23 nsew
rlabel mvndiffc -3870 0 -3870 0 0 S11
port 24 nsew
rlabel polycont -3741 555 -3741 555 0 G11
port 25 nsew
rlabel mvndiffc -3612 0 -3612 0 0 D12
port 26 nsew
rlabel polycont -3483 555 -3483 555 0 G12
port 27 nsew
rlabel mvndiffc -3354 0 -3354 0 0 S13
port 28 nsew
rlabel polycont -3225 555 -3225 555 0 G13
port 29 nsew
rlabel mvndiffc -3096 0 -3096 0 0 D14
port 30 nsew
rlabel polycont -2967 555 -2967 555 0 G14
port 31 nsew
rlabel mvndiffc -2838 0 -2838 0 0 S15
port 32 nsew
rlabel polycont -2709 555 -2709 555 0 G15
port 33 nsew
rlabel mvndiffc -2580 0 -2580 0 0 D16
port 34 nsew
rlabel polycont -2451 555 -2451 555 0 G16
port 35 nsew
rlabel mvndiffc -2322 0 -2322 0 0 S17
port 36 nsew
rlabel polycont -2193 555 -2193 555 0 G17
port 37 nsew
rlabel mvndiffc -2064 0 -2064 0 0 D18
port 38 nsew
rlabel polycont -1935 555 -1935 555 0 G18
port 39 nsew
rlabel mvndiffc -1806 0 -1806 0 0 S19
port 40 nsew
rlabel polycont -1677 555 -1677 555 0 G19
port 41 nsew
rlabel mvndiffc -1548 0 -1548 0 0 D20
port 42 nsew
rlabel polycont -1419 555 -1419 555 0 G20
port 43 nsew
rlabel mvndiffc -1290 0 -1290 0 0 S21
port 44 nsew
rlabel polycont -1161 555 -1161 555 0 G21
port 45 nsew
rlabel mvndiffc -1032 0 -1032 0 0 D22
port 46 nsew
rlabel polycont -903 555 -903 555 0 G22
port 47 nsew
rlabel mvndiffc -774 0 -774 0 0 S23
port 48 nsew
rlabel polycont -645 555 -645 555 0 G23
port 49 nsew
rlabel mvndiffc -516 0 -516 0 0 D24
port 50 nsew
rlabel polycont -387 555 -387 555 0 G24
port 51 nsew
rlabel mvndiffc -258 0 -258 0 0 S25
port 52 nsew
rlabel polycont -129 555 -129 555 0 G25
port 53 nsew
rlabel mvndiffc 0 0 0 0 0 D26
port 54 nsew
rlabel polycont 129 555 129 555 0 G26
port 55 nsew
rlabel mvndiffc 258 0 258 0 0 S27
port 56 nsew
rlabel polycont 387 555 387 555 0 G27
port 57 nsew
rlabel mvndiffc 516 0 516 0 0 D28
port 58 nsew
rlabel polycont 645 555 645 555 0 G28
port 59 nsew
rlabel mvndiffc 774 0 774 0 0 S29
port 60 nsew
rlabel polycont 903 555 903 555 0 G29
port 61 nsew
rlabel mvndiffc 1032 0 1032 0 0 D30
port 62 nsew
rlabel polycont 1161 555 1161 555 0 G30
port 63 nsew
rlabel mvndiffc 1290 0 1290 0 0 S31
port 64 nsew
rlabel polycont 1419 555 1419 555 0 G31
port 65 nsew
rlabel mvndiffc 1548 0 1548 0 0 D32
port 66 nsew
rlabel polycont 1677 555 1677 555 0 G32
port 67 nsew
rlabel mvndiffc 1806 0 1806 0 0 S33
port 68 nsew
rlabel polycont 1935 555 1935 555 0 G33
port 69 nsew
rlabel mvndiffc 2064 0 2064 0 0 D34
port 70 nsew
rlabel polycont 2193 555 2193 555 0 G34
port 71 nsew
rlabel mvndiffc 2322 0 2322 0 0 S35
port 72 nsew
rlabel polycont 2451 555 2451 555 0 G35
port 73 nsew
rlabel mvndiffc 2580 0 2580 0 0 D36
port 74 nsew
rlabel polycont 2709 555 2709 555 0 G36
port 75 nsew
rlabel mvndiffc 2838 0 2838 0 0 S37
port 76 nsew
rlabel polycont 2967 555 2967 555 0 G37
port 77 nsew
rlabel mvndiffc 3096 0 3096 0 0 D38
port 78 nsew
rlabel polycont 3225 555 3225 555 0 G38
port 79 nsew
rlabel mvndiffc 3354 0 3354 0 0 S39
port 80 nsew
rlabel polycont 3483 555 3483 555 0 G39
port 81 nsew
rlabel mvndiffc 3612 0 3612 0 0 D40
port 82 nsew
rlabel polycont 3741 555 3741 555 0 G40
port 83 nsew
rlabel mvndiffc 3870 0 3870 0 0 S41
port 84 nsew
rlabel polycont 3999 555 3999 555 0 G41
port 85 nsew
rlabel mvndiffc 4128 0 4128 0 0 D42
port 86 nsew
rlabel polycont 4257 555 4257 555 0 G42
port 87 nsew
rlabel mvndiffc 4386 0 4386 0 0 S43
port 88 nsew
rlabel polycont 4515 555 4515 555 0 G43
port 89 nsew
rlabel mvndiffc 4644 0 4644 0 0 D44
port 90 nsew
rlabel polycont 4773 555 4773 555 0 G44
port 91 nsew
rlabel mvndiffc 4902 0 4902 0 0 S45
port 92 nsew
rlabel polycont 5031 555 5031 555 0 G45
port 93 nsew
rlabel mvndiffc 5160 0 5160 0 0 D46
port 94 nsew
rlabel polycont 5289 555 5289 555 0 G46
port 95 nsew
rlabel mvndiffc 5418 0 5418 0 0 S47
port 96 nsew
rlabel polycont 5547 555 5547 555 0 G47
port 97 nsew
rlabel mvndiffc 5676 0 5676 0 0 D48
port 98 nsew
rlabel polycont 5805 555 5805 555 0 G48
port 99 nsew
rlabel mvndiffc 5934 0 5934 0 0 S49
port 100 nsew
rlabel polycont 6063 555 6063 555 0 G49
port 101 nsew
rlabel mvndiffc 6192 0 6192 0 0 D50
port 102 nsew
rlabel polycont 6321 555 6321 555 0 G50
port 103 nsew
rlabel mvndiffc 6450 0 6450 0 0 S51
port 104 nsew
rlabel polycont 6579 555 6579 555 0 G51
port 105 nsew
<< properties >>
string FIXED_BBOX -6844 -693 6844 693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 1 m 1 nf 52 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
