magic
tech sky130A
magscale 1 2
timestamp 1756728921
<< viali >>
rect -14 7912 4216 7946
rect -114 6108 -80 7846
rect 4282 6108 4316 7846
rect 4740 7653 7374 7687
rect 4640 6367 4674 7587
rect 7440 6367 7474 7587
rect 4740 6267 7374 6301
rect -14 6008 4216 6042
<< metal1 >>
rect -120 7946 4322 7952
rect -120 7912 -14 7946
rect 4216 7912 4322 7946
rect -120 7906 4322 7912
rect -120 7846 -74 7906
rect -120 7131 -114 7846
rect -123 7125 -114 7131
rect -80 7131 -74 7846
rect 624 7863 740 7869
rect 262 7768 328 7814
rect 882 7863 998 7869
rect 108 7713 224 7719
rect 778 7768 844 7814
rect 1656 7863 1772 7869
rect 366 7713 482 7719
rect 1294 7768 1360 7814
rect 1914 7863 2030 7869
rect 1140 7713 1256 7719
rect 1810 7768 1876 7814
rect 2172 7863 2288 7869
rect 2430 7863 2546 7869
rect 2326 7768 2392 7814
rect 3204 7863 3320 7869
rect 1398 7713 1514 7719
rect 2842 7768 2908 7814
rect 3462 7863 3578 7869
rect 2688 7713 2804 7719
rect 3358 7768 3424 7814
rect 4276 7846 4322 7906
rect 2946 7713 3062 7719
rect 3874 7768 3940 7814
rect 3720 7713 3836 7719
rect 3978 7713 4094 7719
rect 11 7421 63 7427
rect -80 7125 -71 7131
rect -123 6823 -114 6829
rect -120 6108 -114 6823
rect -80 6823 -71 6829
rect -80 6108 -74 6823
rect 11 6527 63 6533
rect 269 7421 321 7427
rect 269 6527 321 6533
rect 527 7421 579 7427
rect 527 6527 579 6533
rect 785 7421 837 7427
rect 785 6527 837 6533
rect 1043 7421 1095 7427
rect 1043 6527 1095 6533
rect 1301 7421 1353 7427
rect 1301 6527 1353 6533
rect 1559 7421 1611 7427
rect 1559 6527 1611 6533
rect 1817 7421 1869 7427
rect 1817 6527 1869 6533
rect 2075 7421 2127 7427
rect 2075 6527 2127 6533
rect 2333 7421 2385 7427
rect 2333 6527 2385 6533
rect 2591 7421 2643 7427
rect 2591 6527 2643 6533
rect 2849 7421 2901 7427
rect 2849 6527 2901 6533
rect 3107 7421 3159 7427
rect 3107 6527 3159 6533
rect 3365 7421 3417 7427
rect 3365 6527 3417 6533
rect 3623 7421 3675 7427
rect 3623 6527 3675 6533
rect 3881 7421 3933 7427
rect 3881 6527 3933 6533
rect 4139 7421 4191 7427
rect 4276 7131 4282 7846
rect 4273 7125 4282 7131
rect 4316 7131 4322 7846
rect 4634 7687 7480 7693
rect 4634 7653 4740 7687
rect 7374 7653 7480 7687
rect 4634 7647 7480 7653
rect 4634 7587 4680 7647
rect 4316 7125 4325 7131
rect 4273 6823 4282 6829
rect 4139 6527 4191 6533
rect 624 6235 740 6241
rect -120 6048 -74 6108
rect 262 6140 328 6186
rect 882 6235 998 6241
rect 108 6085 224 6091
rect 778 6140 844 6186
rect 1656 6235 1772 6241
rect 366 6085 482 6091
rect 1294 6140 1360 6186
rect 1914 6235 2030 6241
rect 1140 6085 1256 6091
rect 1810 6140 1876 6186
rect 2172 6235 2288 6241
rect 2430 6235 2546 6241
rect 2326 6140 2392 6186
rect 3204 6235 3320 6241
rect 1398 6085 1514 6091
rect 2842 6140 2908 6186
rect 3462 6235 3578 6241
rect 2688 6085 2804 6091
rect 3358 6140 3424 6186
rect 2946 6085 3062 6091
rect 3874 6140 3940 6186
rect 3720 6085 3836 6091
rect 3978 6085 4094 6091
rect 4276 6108 4282 6823
rect 4316 6823 4325 6829
rect 4316 6108 4322 6823
rect 4276 6048 4322 6108
rect 4634 6367 4640 7587
rect 4674 6367 4680 7587
rect 4846 7605 4898 7611
rect 5004 7605 5056 7611
rect 4918 7509 4984 7555
rect 5478 7605 5530 7611
rect 5234 7509 5300 7555
rect 5636 7605 5688 7611
rect 5162 7458 5214 7464
rect 5550 7509 5616 7555
rect 6426 7605 6478 7611
rect 5320 7458 5372 7464
rect 5866 7509 5932 7555
rect 5794 7458 5846 7464
rect 5952 7458 6004 7464
rect 6182 7509 6248 7555
rect 6584 7605 6636 7611
rect 6110 7458 6162 7464
rect 6498 7509 6564 7555
rect 7058 7605 7110 7611
rect 6268 7458 6320 7464
rect 6814 7509 6880 7555
rect 7216 7605 7268 7611
rect 6742 7458 6794 7464
rect 7130 7509 7196 7555
rect 7434 7587 7480 7647
rect 6900 7458 6952 7464
rect 4767 7421 4819 7427
rect 4767 6527 4819 6533
rect 4925 7421 4977 7427
rect 4925 6527 4977 6533
rect 5083 7421 5135 7427
rect 5083 6527 5135 6533
rect 5241 7421 5293 7427
rect 5241 6527 5293 6533
rect 5399 7421 5451 7427
rect 5399 6527 5451 6533
rect 5557 7421 5609 7427
rect 5557 6527 5609 6533
rect 5715 7421 5767 7427
rect 5715 6527 5767 6533
rect 5873 7421 5925 7427
rect 5873 6527 5925 6533
rect 6031 7421 6083 7427
rect 6031 6527 6083 6533
rect 6189 7421 6241 7427
rect 6189 6527 6241 6533
rect 6347 7421 6399 7427
rect 6347 6527 6399 6533
rect 6505 7421 6557 7427
rect 6505 6527 6557 6533
rect 6663 7421 6715 7427
rect 6663 6527 6715 6533
rect 6821 7421 6873 7427
rect 6821 6527 6873 6533
rect 6979 7421 7031 7427
rect 6979 6527 7031 6533
rect 7137 7421 7189 7427
rect 7137 6527 7189 6533
rect 7295 7421 7347 7427
rect 7295 6527 7347 6533
rect 4846 6490 4898 6496
rect 5004 6490 5056 6496
rect 4918 6399 4984 6445
rect 5478 6490 5530 6496
rect 4634 6307 4680 6367
rect 5234 6399 5300 6445
rect 5636 6490 5688 6496
rect 5162 6343 5214 6349
rect 5550 6399 5616 6445
rect 6426 6490 6478 6496
rect 5320 6343 5372 6349
rect 5866 6399 5932 6445
rect 5794 6343 5846 6349
rect 5952 6343 6004 6349
rect 6182 6399 6248 6445
rect 6584 6490 6636 6496
rect 6110 6343 6162 6349
rect 6498 6399 6564 6445
rect 7058 6490 7110 6496
rect 6268 6343 6320 6349
rect 6814 6399 6880 6445
rect 7216 6490 7268 6496
rect 6742 6343 6794 6349
rect 7130 6399 7196 6445
rect 6900 6343 6952 6349
rect 7434 6367 7440 7587
rect 7474 6367 7480 7587
rect 7434 6307 7480 6367
rect 4634 6301 7480 6307
rect 7374 6267 7480 6301
rect 4770 6261 7480 6267
rect 4634 6077 4770 6083
rect -120 6042 4322 6048
rect -120 6008 -14 6042
rect 4216 6008 4322 6042
rect -120 6002 4322 6008
<< via1 >>
rect 108 7719 224 7771
rect 624 7811 740 7863
rect 366 7719 482 7771
rect 882 7811 998 7863
rect 1140 7719 1256 7771
rect 1656 7811 1772 7863
rect 1398 7719 1514 7771
rect 1914 7811 2030 7863
rect 2172 7811 2288 7863
rect 2430 7811 2546 7863
rect 2688 7719 2804 7771
rect 3204 7811 3320 7863
rect 2946 7719 3062 7771
rect 3462 7811 3578 7863
rect 3720 7719 3836 7771
rect 3978 7719 4094 7771
rect -123 6829 -114 7125
rect -114 6829 -80 7125
rect -80 6829 -71 7125
rect 11 6533 63 7421
rect 269 6533 321 7421
rect 527 6533 579 7421
rect 785 6533 837 7421
rect 1043 6533 1095 7421
rect 1301 6533 1353 7421
rect 1559 6533 1611 7421
rect 1817 6533 1869 7421
rect 2075 6533 2127 7421
rect 2333 6533 2385 7421
rect 2591 6533 2643 7421
rect 2849 6533 2901 7421
rect 3107 6533 3159 7421
rect 3365 6533 3417 7421
rect 3623 6533 3675 7421
rect 3881 6533 3933 7421
rect 4139 6533 4191 7421
rect 4273 6829 4282 7125
rect 4282 6829 4316 7125
rect 4316 6829 4325 7125
rect 108 6091 224 6143
rect 624 6183 740 6235
rect 366 6091 482 6143
rect 882 6183 998 6235
rect 1140 6091 1256 6143
rect 1656 6183 1772 6235
rect 1398 6091 1514 6143
rect 1914 6183 2030 6235
rect 2172 6183 2288 6235
rect 2430 6183 2546 6235
rect 2688 6091 2804 6143
rect 3204 6183 3320 6235
rect 2946 6091 3062 6143
rect 3462 6183 3578 6235
rect 3720 6091 3836 6143
rect 3978 6091 4094 6143
rect 4846 7553 4898 7605
rect 5004 7553 5056 7605
rect 5162 7464 5214 7516
rect 5478 7553 5530 7605
rect 5320 7464 5372 7516
rect 5636 7553 5688 7605
rect 5794 7464 5846 7516
rect 5952 7464 6004 7516
rect 6110 7464 6162 7516
rect 6426 7553 6478 7605
rect 6268 7464 6320 7516
rect 6584 7553 6636 7605
rect 6742 7464 6794 7516
rect 7058 7553 7110 7605
rect 6900 7464 6952 7516
rect 7216 7553 7268 7605
rect 4767 6533 4819 7421
rect 4925 6533 4977 7421
rect 5083 6533 5135 7421
rect 5241 6533 5293 7421
rect 5399 6533 5451 7421
rect 5557 6533 5609 7421
rect 5715 6533 5767 7421
rect 5873 6533 5925 7421
rect 6031 6533 6083 7421
rect 6189 6533 6241 7421
rect 6347 6533 6399 7421
rect 6505 6533 6557 7421
rect 6663 6533 6715 7421
rect 6821 6533 6873 7421
rect 6979 6533 7031 7421
rect 7137 6533 7189 7421
rect 7295 6533 7347 7421
rect 4846 6438 4898 6490
rect 5004 6438 5056 6490
rect 5162 6349 5214 6401
rect 5478 6438 5530 6490
rect 5320 6349 5372 6401
rect 5636 6438 5688 6490
rect 5794 6349 5846 6401
rect 5952 6349 6004 6401
rect 6110 6349 6162 6401
rect 6426 6438 6478 6490
rect 6268 6349 6320 6401
rect 6584 6438 6636 6490
rect 6742 6349 6794 6401
rect 7058 6438 7110 6490
rect 6900 6349 6952 6401
rect 7216 6438 7268 6490
rect 4634 6267 4740 6301
rect 4740 6267 4770 6301
rect 4634 6083 4770 6267
<< metal2 >>
rect 1640 8051 1940 8056
rect 1640 7863 1649 8051
rect 1931 7863 1940 8051
rect 70 7811 624 7863
rect 740 7811 882 7863
rect 998 7861 1649 7863
rect 998 7811 1656 7861
rect 1772 7811 1914 7861
rect 2030 7811 2172 7863
rect 2288 7811 2430 7863
rect 2546 7811 3204 7863
rect 3320 7811 3462 7863
rect 3578 7811 4431 7863
rect -229 7719 108 7771
rect 224 7719 366 7771
rect 482 7719 1140 7771
rect 1256 7719 1398 7771
rect 1514 7719 2688 7771
rect 2804 7719 2946 7771
rect 3062 7719 3720 7771
rect 3836 7719 3978 7771
rect 4094 7719 4132 7771
rect -229 6143 -177 7719
rect 11 7421 63 7427
rect -125 7125 -69 7131
rect -125 7122 -123 7125
rect -71 7122 -69 7125
rect -125 6829 -123 6832
rect -71 6829 -69 6832
rect -125 6823 -69 6829
rect 9 7122 11 7131
rect 269 7421 321 7427
rect 63 7122 65 7131
rect 9 6823 11 6832
rect 63 6823 65 6832
rect 11 6527 63 6533
rect 227 6718 269 6727
rect 527 7421 579 7427
rect 485 7122 527 7131
rect 743 7421 879 7427
rect 743 7418 785 7421
rect 837 7418 879 7421
rect 743 7227 785 7236
rect 579 7122 621 7131
rect 485 6823 527 6832
rect 321 6718 363 6727
rect 227 6533 269 6536
rect 321 6533 363 6536
rect 227 6527 363 6533
rect 579 6823 621 6832
rect 527 6527 579 6533
rect 837 7227 879 7236
rect 1043 7421 1095 7427
rect 1001 7122 1043 7131
rect 1301 7421 1353 7427
rect 1095 7122 1137 7131
rect 1001 6823 1043 6832
rect 785 6527 837 6533
rect 1095 6823 1137 6832
rect 1043 6527 1095 6533
rect 1259 6718 1301 6727
rect 1559 7421 1611 7427
rect 1517 7122 1559 7131
rect 1775 7421 1911 7427
rect 1775 7418 1817 7421
rect 1869 7418 1911 7421
rect 1775 7227 1817 7236
rect 1611 7122 1653 7131
rect 1517 6823 1559 6832
rect 1353 6718 1395 6727
rect 1259 6533 1301 6536
rect 1353 6533 1395 6536
rect 1259 6527 1395 6533
rect 1611 6823 1653 6832
rect 1559 6527 1611 6533
rect 1869 7227 1911 7236
rect 2075 7421 2127 7427
rect 2033 7122 2075 7131
rect 2291 7421 2427 7427
rect 2291 7418 2333 7421
rect 2385 7418 2427 7421
rect 2291 7227 2333 7236
rect 2127 7122 2169 7131
rect 2033 6823 2075 6832
rect 1817 6527 1869 6533
rect 2127 6823 2169 6832
rect 2075 6527 2127 6533
rect 2385 7227 2427 7236
rect 2591 7421 2643 7427
rect 2549 7122 2591 7131
rect 2849 7421 2901 7427
rect 2643 7122 2685 7131
rect 2549 6823 2591 6832
rect 2333 6527 2385 6533
rect 2643 6823 2685 6832
rect 2591 6527 2643 6533
rect 2807 6718 2849 6727
rect 3107 7421 3159 7427
rect 3065 7122 3107 7131
rect 3323 7421 3459 7427
rect 3323 7418 3365 7421
rect 3417 7418 3459 7421
rect 3323 7227 3365 7236
rect 3159 7122 3201 7131
rect 3065 6823 3107 6832
rect 2901 6718 2943 6727
rect 2807 6533 2849 6536
rect 2901 6533 2943 6536
rect 2807 6527 2943 6533
rect 3159 6823 3201 6832
rect 3107 6527 3159 6533
rect 3417 7227 3459 7236
rect 3623 7421 3675 7427
rect 3581 7122 3623 7131
rect 3881 7421 3933 7427
rect 3675 7122 3717 7131
rect 3581 6823 3623 6832
rect 3365 6527 3417 6533
rect 3675 6823 3717 6832
rect 3623 6527 3675 6533
rect 3839 6718 3881 6727
rect 4139 7421 4191 7427
rect 4137 7122 4139 7131
rect 4191 7122 4193 7131
rect 4137 6823 4139 6832
rect 3933 6718 3975 6727
rect 3839 6533 3881 6536
rect 3933 6533 3975 6536
rect 3839 6527 3975 6533
rect 4191 6823 4193 6832
rect 4271 7125 4327 7131
rect 4271 7122 4273 7125
rect 4325 7122 4327 7125
rect 4271 6829 4273 6832
rect 4325 6829 4327 6832
rect 4271 6823 4327 6829
rect 4139 6527 4191 6533
rect 4379 6235 4431 7811
rect 4485 7744 4631 7753
rect 4485 7562 4490 7744
rect 4626 7605 4631 7744
rect 7483 7655 7629 7664
rect 4626 7562 4846 7605
rect 4485 7553 4846 7562
rect 4898 7553 5004 7605
rect 5056 7553 5478 7605
rect 5530 7553 5636 7605
rect 5688 7553 6426 7605
rect 6478 7553 6584 7605
rect 6636 7553 7058 7605
rect 7110 7553 7216 7605
rect 7268 7553 7288 7605
rect 4631 6490 4683 7553
rect 7483 7516 7488 7655
rect 4826 7464 5162 7516
rect 5214 7464 5320 7516
rect 5372 7464 5794 7516
rect 5846 7464 5952 7516
rect 6004 7464 6110 7516
rect 6162 7464 6268 7516
rect 6320 7464 6742 7516
rect 6794 7464 6900 7516
rect 6952 7473 7488 7516
rect 7624 7473 7629 7655
rect 6952 7464 7629 7473
rect 4767 7421 4819 7427
rect 4765 7122 4767 7131
rect 4883 7421 5019 7427
rect 4883 7418 4925 7421
rect 4977 7418 5019 7421
rect 4883 7227 4925 7236
rect 4819 7122 4821 7131
rect 4765 6823 4767 6832
rect 4819 6823 4821 6832
rect 4767 6527 4819 6533
rect 4977 7227 5019 7236
rect 5083 7421 5135 7427
rect 5041 7122 5083 7131
rect 5241 7421 5293 7427
rect 5135 7122 5177 7131
rect 5041 6823 5083 6832
rect 4925 6527 4977 6533
rect 5135 6823 5177 6832
rect 5083 6527 5135 6533
rect 5199 6718 5241 6727
rect 5399 7421 5451 7427
rect 5357 7122 5399 7131
rect 5515 7421 5651 7427
rect 5515 7418 5557 7421
rect 5609 7418 5651 7421
rect 5515 7227 5557 7236
rect 5451 7122 5493 7131
rect 5357 6823 5399 6832
rect 5293 6718 5335 6727
rect 5199 6533 5241 6536
rect 5293 6533 5335 6536
rect 5199 6527 5335 6533
rect 5451 6823 5493 6832
rect 5399 6527 5451 6533
rect 5609 7227 5651 7236
rect 5715 7421 5767 7427
rect 5673 7122 5715 7131
rect 5873 7421 5925 7427
rect 5767 7122 5809 7131
rect 5673 6823 5715 6832
rect 5557 6527 5609 6533
rect 5767 6823 5809 6832
rect 5715 6527 5767 6533
rect 5831 6718 5873 6727
rect 6031 7421 6083 7427
rect 5989 7122 6031 7131
rect 6189 7421 6241 7427
rect 6083 7122 6125 7131
rect 5989 6823 6031 6832
rect 5925 6718 5967 6727
rect 5831 6533 5873 6536
rect 5925 6533 5967 6536
rect 5831 6527 5967 6533
rect 6083 6823 6125 6832
rect 6031 6527 6083 6533
rect 6147 6718 6189 6727
rect 6347 7421 6399 7427
rect 6305 7122 6347 7131
rect 6463 7421 6599 7427
rect 6463 7418 6505 7421
rect 6557 7418 6599 7421
rect 6463 7227 6505 7236
rect 6399 7122 6441 7131
rect 6305 6823 6347 6832
rect 6241 6718 6283 6727
rect 6147 6533 6189 6536
rect 6241 6533 6283 6536
rect 6147 6527 6283 6533
rect 6399 6823 6441 6832
rect 6347 6527 6399 6533
rect 6557 7227 6599 7236
rect 6663 7421 6715 7427
rect 6621 7122 6663 7131
rect 6821 7421 6873 7427
rect 6715 7122 6757 7131
rect 6621 6823 6663 6832
rect 6505 6527 6557 6533
rect 6715 6823 6757 6832
rect 6663 6527 6715 6533
rect 6779 6718 6821 6727
rect 6979 7421 7031 7427
rect 6937 7122 6979 7131
rect 7095 7421 7231 7427
rect 7095 7418 7137 7421
rect 7189 7418 7231 7421
rect 7095 7227 7137 7236
rect 7031 7122 7073 7131
rect 6937 6823 6979 6832
rect 6873 6718 6915 6727
rect 6779 6533 6821 6536
rect 6873 6533 6915 6536
rect 6779 6527 6915 6533
rect 7031 6823 7073 6832
rect 6979 6527 7031 6533
rect 7189 7227 7231 7236
rect 7295 7421 7347 7427
rect 7293 7122 7295 7131
rect 7347 7122 7349 7131
rect 7293 6823 7295 6832
rect 7137 6527 7189 6533
rect 7347 6823 7349 6832
rect 7295 6527 7347 6533
rect 4631 6438 4846 6490
rect 4898 6438 5004 6490
rect 5056 6438 5478 6490
rect 5530 6438 5636 6490
rect 5688 6438 6426 6490
rect 6478 6438 6584 6490
rect 6636 6438 7058 6490
rect 7110 6438 7216 6490
rect 7268 6438 7288 6490
rect 7431 6401 7483 7464
rect 4826 6349 5162 6401
rect 5214 6349 5320 6401
rect 5372 6349 5794 6401
rect 5846 6349 5952 6401
rect 6004 6349 6110 6401
rect 6162 6349 6268 6401
rect 6320 6349 6742 6401
rect 6794 6349 6900 6401
rect 6952 6349 7483 6401
rect 70 6183 624 6235
rect 740 6183 882 6235
rect 998 6183 1656 6235
rect 1772 6183 1914 6235
rect 2030 6183 2172 6235
rect 2288 6183 2430 6235
rect 2546 6183 3204 6235
rect 3320 6183 3462 6235
rect 3578 6183 4431 6235
rect 4634 6301 4770 6307
rect -229 6091 108 6143
rect 224 6091 366 6143
rect 482 6091 1140 6143
rect 1256 6091 1398 6143
rect 1514 6093 2688 6143
rect 1514 6091 1649 6093
rect 1640 5903 1649 6091
rect 1931 6091 2688 6093
rect 2804 6091 2946 6143
rect 3062 6091 3720 6143
rect 3836 6091 3978 6143
rect 4094 6091 4132 6143
rect 1931 5903 1940 6091
rect 4634 6077 4770 6083
rect 1640 5898 1940 5903
<< via2 >>
rect 1649 7863 1931 8051
rect 1649 7861 1656 7863
rect 1656 7861 1772 7863
rect 1772 7861 1914 7863
rect 1914 7861 1931 7863
rect -125 6832 -123 7122
rect -123 6832 -71 7122
rect -71 6832 -69 7122
rect 9 6832 11 7122
rect 11 6832 63 7122
rect 63 6832 65 7122
rect 743 7236 785 7418
rect 785 7236 837 7418
rect 837 7236 879 7418
rect 485 6832 527 7122
rect 527 6832 579 7122
rect 579 6832 621 7122
rect 227 6536 269 6718
rect 269 6536 321 6718
rect 321 6536 363 6718
rect 1001 6832 1043 7122
rect 1043 6832 1095 7122
rect 1095 6832 1137 7122
rect 1775 7236 1817 7418
rect 1817 7236 1869 7418
rect 1869 7236 1911 7418
rect 1517 6832 1559 7122
rect 1559 6832 1611 7122
rect 1611 6832 1653 7122
rect 1259 6536 1301 6718
rect 1301 6536 1353 6718
rect 1353 6536 1395 6718
rect 2291 7236 2333 7418
rect 2333 7236 2385 7418
rect 2385 7236 2427 7418
rect 2033 6832 2075 7122
rect 2075 6832 2127 7122
rect 2127 6832 2169 7122
rect 2549 6832 2591 7122
rect 2591 6832 2643 7122
rect 2643 6832 2685 7122
rect 3323 7236 3365 7418
rect 3365 7236 3417 7418
rect 3417 7236 3459 7418
rect 3065 6832 3107 7122
rect 3107 6832 3159 7122
rect 3159 6832 3201 7122
rect 2807 6536 2849 6718
rect 2849 6536 2901 6718
rect 2901 6536 2943 6718
rect 3581 6832 3623 7122
rect 3623 6832 3675 7122
rect 3675 6832 3717 7122
rect 4137 6832 4139 7122
rect 4139 6832 4191 7122
rect 4191 6832 4193 7122
rect 3839 6536 3881 6718
rect 3881 6536 3933 6718
rect 3933 6536 3975 6718
rect 4271 6832 4273 7122
rect 4273 6832 4325 7122
rect 4325 6832 4327 7122
rect 4490 7562 4626 7744
rect 7488 7473 7624 7655
rect 4883 7236 4925 7418
rect 4925 7236 4977 7418
rect 4977 7236 5019 7418
rect 4765 6832 4767 7122
rect 4767 6832 4819 7122
rect 4819 6832 4821 7122
rect 5041 6832 5083 7122
rect 5083 6832 5135 7122
rect 5135 6832 5177 7122
rect 5515 7236 5557 7418
rect 5557 7236 5609 7418
rect 5609 7236 5651 7418
rect 5357 6832 5399 7122
rect 5399 6832 5451 7122
rect 5451 6832 5493 7122
rect 5199 6536 5241 6718
rect 5241 6536 5293 6718
rect 5293 6536 5335 6718
rect 5673 6832 5715 7122
rect 5715 6832 5767 7122
rect 5767 6832 5809 7122
rect 5989 6832 6031 7122
rect 6031 6832 6083 7122
rect 6083 6832 6125 7122
rect 5831 6536 5873 6718
rect 5873 6536 5925 6718
rect 5925 6536 5967 6718
rect 6463 7236 6505 7418
rect 6505 7236 6557 7418
rect 6557 7236 6599 7418
rect 6305 6832 6347 7122
rect 6347 6832 6399 7122
rect 6399 6832 6441 7122
rect 6147 6536 6189 6718
rect 6189 6536 6241 6718
rect 6241 6536 6283 6718
rect 6621 6832 6663 7122
rect 6663 6832 6715 7122
rect 6715 6832 6757 7122
rect 7095 7236 7137 7418
rect 7137 7236 7189 7418
rect 7189 7236 7231 7418
rect 6937 6832 6979 7122
rect 6979 6832 7031 7122
rect 7031 6832 7073 7122
rect 6779 6536 6821 6718
rect 6821 6536 6873 6718
rect 6873 6536 6915 6718
rect 7293 6832 7295 7122
rect 7295 6832 7347 7122
rect 7347 6832 7349 7122
rect 1649 5903 1931 6093
rect 4634 6086 4770 6268
<< metal3 >>
rect 5970 12897 6270 12898
rect 5970 12699 5976 12897
rect 6264 12699 6270 12897
rect 5970 12698 6270 12699
rect 6570 12897 6870 12898
rect 6570 12699 6576 12897
rect 6864 12699 6870 12897
rect 6570 12698 6870 12699
rect 1644 8051 1936 8056
rect 1644 7861 1649 8051
rect 1931 7861 1936 8051
rect 6047 8049 6193 12698
rect 1644 7427 1936 7861
rect 4485 7903 6193 8049
rect 6647 8049 6793 12698
rect 6647 7903 7629 8049
rect 4485 7744 4631 7903
rect 4485 7562 4490 7744
rect 4626 7562 4631 7744
rect 4485 7553 4631 7562
rect 7483 7655 7629 7903
rect 7483 7473 7488 7655
rect 7624 7473 7629 7655
rect 7483 7464 7629 7473
rect -1390 7426 7236 7427
rect -1390 7228 -1384 7426
rect -1096 7418 5971 7426
rect -1096 7236 743 7418
rect 879 7236 1775 7418
rect 1911 7236 2291 7418
rect 2427 7236 3323 7418
rect 3459 7236 4883 7418
rect 5019 7236 5515 7418
rect 5651 7236 5971 7418
rect -1096 7228 5971 7236
rect 6269 7418 7236 7426
rect 6269 7236 6463 7418
rect 6599 7236 7095 7418
rect 7231 7236 7236 7418
rect 6269 7228 7236 7236
rect -1390 7227 7236 7228
rect -140 7126 4332 7127
rect -140 7122 666 7126
rect -140 6832 -125 7122
rect -69 6832 9 7122
rect 65 6832 485 7122
rect 621 6832 666 7122
rect -140 6828 666 6832
rect 894 7122 4332 7126
rect 894 6832 1001 7122
rect 1137 6832 1517 7122
rect 1653 6832 2033 7122
rect 2169 6832 2549 7122
rect 2685 6832 3065 7122
rect 3201 6832 3581 7122
rect 3717 6832 4137 7122
rect 4193 6832 4271 7122
rect 4327 6832 4332 7122
rect 894 6828 4332 6832
rect -140 6827 4332 6828
rect 4760 7122 7354 7127
rect 4760 6832 4765 7122
rect 4821 6832 5041 7122
rect 5177 6832 5357 7122
rect 5493 6832 5673 7122
rect 5809 6832 5989 7122
rect 6125 6832 6305 7122
rect 6441 6832 6621 7122
rect 6757 6832 6937 7122
rect 7073 6832 7293 7122
rect 7349 6832 7354 7122
rect 4760 6827 7354 6832
rect -78 6726 6920 6727
rect -78 6718 2296 6726
rect -78 6536 227 6718
rect 363 6536 1259 6718
rect 1395 6536 2296 6718
rect -78 6528 2296 6536
rect 2584 6718 6920 6726
rect 2584 6536 2807 6718
rect 2943 6536 3839 6718
rect 3975 6536 5199 6718
rect 5335 6536 5831 6718
rect 5967 6536 6147 6718
rect 6283 6536 6779 6718
rect 6915 6536 6920 6718
rect 2584 6528 6920 6536
rect -78 6527 6920 6528
rect 4020 6276 4775 6277
rect 1640 6093 1940 6098
rect 1640 5903 1649 6093
rect 1931 5903 1940 6093
rect 4020 6078 4026 6276
rect 4254 6268 4775 6276
rect 4254 6086 4634 6268
rect 4770 6086 4775 6268
rect 4254 6078 4775 6086
rect 4020 6077 4775 6078
rect 1640 4262 1940 5903
rect 1640 3962 3980 4262
rect 1640 3628 1940 3962
rect 3680 3628 3980 3962
rect 954 1224 1001 1288
rect 1065 1224 1071 1288
rect 4634 1224 4681 1288
rect 4745 1224 4751 1288
<< via3 >>
rect 5976 12699 6264 12897
rect 6576 12699 6864 12897
rect -1384 7228 -1096 7426
rect 5971 7228 6269 7426
rect 666 6828 894 7126
rect 2296 6528 2584 6726
rect 4026 6078 4254 6276
rect 2291 1525 2589 1923
rect 5971 1525 6269 1923
rect 1001 1224 1065 1288
rect 4681 1224 4745 1288
<< metal4 >>
rect -1390 7426 -1090 12998
rect -1390 7228 -1384 7426
rect -1096 7228 -1090 7426
rect -1390 7227 -1090 7228
rect 20 5576 260 12998
rect 340 5576 580 12998
rect 660 7126 900 12998
rect 660 6828 666 7126
rect 894 6828 900 7126
rect 660 5576 900 6828
rect 2290 6726 2590 12998
rect 2290 6528 2296 6726
rect 2584 6528 2590 6726
rect 2290 1923 2590 6528
rect 3700 5576 3940 12998
rect 4020 6276 4260 12998
rect 4020 6078 4026 6276
rect 4254 6078 4260 6276
rect 4020 5576 4260 6078
rect 4340 5576 4580 12998
rect 5970 12897 6270 12998
rect 5970 12699 5976 12897
rect 6264 12699 6270 12897
rect 5970 12698 6270 12699
rect 6570 12897 6870 12998
rect 6570 12699 6576 12897
rect 6864 12699 6870 12897
rect 6570 12698 6870 12699
rect 5970 7426 6270 7427
rect 5970 7228 5971 7426
rect 6269 7228 6270 7426
rect 2290 1525 2291 1923
rect 2589 1525 2590 1923
rect 2290 1524 2590 1525
rect 5970 1923 6270 7228
rect 5970 1525 5971 1923
rect 6269 1525 6270 1923
rect 5970 1524 6270 1525
rect 1000 1288 1066 1289
rect 1000 1224 1001 1288
rect 1065 1224 1066 1288
rect 4680 1288 4746 1289
rect 4680 1224 4681 1288
rect 4745 1224 4746 1288
rect 20 1136 260 1224
rect 340 1136 580 1224
rect 660 -48 900 1224
rect 1000 1221 1066 1224
rect 1000 1140 1060 1221
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1221 4746 1224
rect 4680 1140 4740 1221
use dev_ctrl_b1  dev_ctrl_b1_0
timestamp 1756101716
transform 1 0 3680 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e1  dev_ctrl_e1_0
timestamp 1756101705
transform 1 0 0 0 1 0
box -38 -48 6868 1140
use sky130_fd_pr__nfet_g5v0d10v5_WZKDHM  sky130_fd_pr__nfet_g5v0d10v5_WZKDHM_0
timestamp 1756220169
transform 1 0 6057 0 1 6977
box -1465 -758 1465 758
use sky130_fd_pr__pfet_g5v0d10v5_L2ZWMC  sky130_fd_pr__pfet_g5v0d10v5_L2ZWMC_0
timestamp 1756728921
transform 1 0 2101 0 1 6977
box -2293 -1047 2293 1047
use tt_asw_3v3  tt_asw_3v3_0
array 0 1 3680 0 0 -4352
timestamp 1756064685
transform 1 0 0 0 -1 5576
box 0 0 3680 4352
<< end >>
