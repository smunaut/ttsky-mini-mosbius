magic
tech sky130A
magscale 1 2
timestamp 1756064830
<< viali >>
rect 1777 833 1811 867
rect 3617 833 3651 867
rect 1501 765 1535 799
rect 3341 765 3375 799
rect 29 629 63 663
rect 1869 629 1903 663
rect 121 425 155 459
rect 949 289 983 323
rect 1501 289 1535 323
rect 765 221 799 255
rect 1133 221 1167 255
rect 1317 221 1351 255
rect 1685 221 1719 255
rect 1869 221 1903 255
<< metal1 >>
rect 1854 960 1860 1012
rect 1912 1000 1918 1012
rect 3694 1000 3700 1012
rect 1912 972 3700 1000
rect 1912 960 1918 972
rect 3694 960 3700 972
rect 3752 1000 3758 1012
rect 3752 972 6868 1000
rect 3752 960 3758 972
rect 400 904 5948 932
rect 1765 867 1823 873
rect 1765 833 1777 867
rect 1811 864 1823 867
rect 1854 864 1860 876
rect 1811 836 1860 864
rect 1811 833 1823 836
rect 1765 827 1823 833
rect 1854 824 1860 836
rect 1912 824 1918 876
rect 3605 867 3663 873
rect 3605 833 3617 867
rect 3651 864 3663 867
rect 3694 864 3700 876
rect 3651 836 3700 864
rect 3651 833 3663 836
rect 3605 827 3663 833
rect 3694 824 3700 836
rect 3752 824 3758 876
rect 1489 799 1547 805
rect 1489 765 1501 799
rect 1535 796 1547 799
rect 1535 768 1716 796
rect 1535 765 1547 768
rect 1489 759 1547 765
rect 17 663 75 669
rect 17 629 29 663
rect 63 660 75 663
rect 1302 660 1308 672
rect 63 632 1308 660
rect 63 629 75 632
rect 17 623 75 629
rect 1302 620 1308 632
rect 1360 620 1366 672
rect 1688 660 1716 768
rect 3326 756 3332 808
rect 3384 756 3390 808
rect 1854 660 1860 672
rect 1688 632 1860 660
rect 1854 620 1860 632
rect 1912 620 1918 672
rect 109 459 167 465
rect 109 456 121 459
rect 32 428 121 456
rect 109 425 121 428
rect 155 425 167 459
rect 109 419 167 425
rect 768 428 1348 456
rect 768 267 796 428
rect 934 280 940 332
rect 992 280 998 332
rect 759 255 805 267
rect 759 221 765 255
rect 799 221 805 255
rect 759 209 805 221
rect 1127 255 1173 267
rect 1320 264 1348 428
rect 3326 416 3332 468
rect 3384 456 3390 468
rect 3384 428 3740 456
rect 3384 416 3390 428
rect 1486 280 1492 332
rect 1544 280 1550 332
rect 1127 221 1133 255
rect 1167 221 1173 255
rect 1127 209 1173 221
rect 1302 212 1308 264
rect 1360 212 1366 264
rect 1679 255 1725 267
rect 1679 221 1685 255
rect 1719 221 1725 255
rect 1679 209 1725 221
rect 1854 212 1860 264
rect 1912 212 1918 264
rect 1136 116 1164 209
rect 1688 116 1716 209
rect 1136 88 5396 116
<< via1 >>
rect 340 1046 580 1130
rect 1860 960 1912 1012
rect 3700 960 3752 1012
rect 1860 824 1912 876
rect 3700 824 3752 876
rect 1308 620 1360 672
rect 3332 799 3384 808
rect 3332 765 3341 799
rect 3341 765 3375 799
rect 3375 765 3384 799
rect 3332 756 3384 765
rect 1860 663 1912 672
rect 1860 629 1869 663
rect 1869 629 1903 663
rect 1903 629 1912 663
rect 1860 620 1912 629
rect 20 502 260 586
rect 940 323 992 332
rect 940 289 949 323
rect 949 289 983 323
rect 983 289 992 323
rect 940 280 992 289
rect 3332 416 3384 468
rect 1492 323 1544 332
rect 1492 289 1501 323
rect 1501 289 1535 323
rect 1535 289 1544 323
rect 1492 280 1544 289
rect 1308 255 1360 264
rect 1308 221 1317 255
rect 1317 221 1351 255
rect 1351 221 1360 255
rect 1308 212 1360 221
rect 1860 255 1912 264
rect 1860 221 1869 255
rect 1869 221 1903 255
rect 1903 221 1912 255
rect 1860 212 1912 221
rect 340 -42 580 42
<< metal2 >>
rect 340 1130 580 1136
rect 340 1040 580 1046
rect 1860 1012 1912 1018
rect 1860 954 1912 960
rect 3700 1012 3752 1018
rect 3700 954 3752 960
rect 1872 882 1900 954
rect 3712 882 3740 954
rect 1860 876 1912 882
rect 938 810 994 819
rect 938 745 994 754
rect 1490 810 1546 819
rect 1860 818 1912 824
rect 3700 876 3752 882
rect 3700 818 3752 824
rect 1490 745 1546 754
rect 3332 808 3384 814
rect 3332 750 3384 756
rect 20 586 260 592
rect 20 496 260 502
rect 952 338 980 745
rect 1308 672 1360 678
rect 1308 614 1360 620
rect 940 332 992 338
rect 940 274 992 280
rect 1320 270 1348 614
rect 1504 338 1532 745
rect 1860 672 1912 678
rect 1860 614 1912 620
rect 1492 332 1544 338
rect 1492 274 1544 280
rect 1872 270 1900 614
rect 3344 474 3372 750
rect 3332 468 3384 474
rect 3332 410 3384 416
rect 1308 264 1360 270
rect 1308 206 1360 212
rect 1860 264 1912 270
rect 1860 206 1912 212
rect 340 42 580 48
rect 340 -48 580 -42
<< via2 >>
rect 345 1049 575 1127
rect 938 754 994 810
rect 1490 754 1546 810
rect 25 505 255 583
rect 345 -39 575 39
<< metal3 >>
rect 340 1130 580 1136
rect 340 1046 341 1130
rect 579 1046 580 1130
rect 340 1040 580 1046
rect 933 814 1060 820
rect 933 810 995 814
rect 933 754 938 810
rect 994 754 995 810
rect 933 750 995 754
rect 1059 750 1060 814
rect 933 744 1060 750
rect 1120 814 1551 820
rect 1120 750 1121 814
rect 1185 810 1551 814
rect 1185 754 1490 810
rect 1546 754 1551 810
rect 1185 750 1551 754
rect 1120 744 1551 750
rect 20 586 260 592
rect 20 502 21 586
rect 259 502 260 586
rect 20 496 260 502
rect 0 372 3680 432
rect 0 242 3680 302
rect 0 112 3680 172
rect 340 42 580 48
rect 340 -42 341 42
rect 579 -42 580 42
rect 340 -48 580 -42
<< via3 >>
rect 341 1127 579 1130
rect 341 1049 345 1127
rect 345 1049 575 1127
rect 575 1049 579 1127
rect 341 1046 579 1049
rect 995 750 1059 814
rect 1121 750 1185 814
rect 21 583 259 586
rect 21 505 25 583
rect 25 505 255 583
rect 255 505 259 583
rect 21 502 259 505
rect 341 39 579 42
rect 341 -39 345 39
rect 345 -39 575 39
rect 575 -39 579 39
rect 341 -42 579 -39
<< metal4 >>
rect 20 586 260 1136
rect 20 502 21 586
rect 259 502 260 586
rect 20 -48 260 502
rect 340 1130 580 1136
rect 340 1046 341 1130
rect 579 1046 580 1130
rect 340 42 580 1046
rect 1000 815 1060 1140
rect 994 814 1060 815
rect 994 750 995 814
rect 1059 750 1060 814
rect 994 749 1060 750
rect 1120 815 1180 1140
rect 1120 814 1186 815
rect 1120 750 1121 814
rect 1185 750 1186 814
rect 1120 749 1186 750
rect 340 -42 341 42
rect 579 -42 580 42
rect 340 -48 580 -42
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform -1 0 1380 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  sky130_fd_sc_hd__and2_2_1
timestamp 1755005639
transform -1 0 1932 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s50_2  sky130_fd_sc_hd__clkdlybuf4s50_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform -1 0 828 0 1 0
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 3128 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 2024 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform -1 0 1840 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sky130_fd_sc_hd__dfrtp_1_1
timestamp 1755005639
transform -1 0 3680 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 3496 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 1932 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755005639
transform 1 0 3588 0 1 0
box -38 -48 130 592
<< labels >>
flabel metal4 20 -48 260 1136 1 FreeSans 160 0 0 0 VDPWR
port 1 n power input
flabel metal4 340 -48 580 1136 1 FreeSans 160 0 0 0 VGND
port 0 n ground input
<< properties >>
string FIXED_BBOX 0 0 3680 1088
<< end >>
