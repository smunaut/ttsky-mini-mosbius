magic
tech sky130A
magscale 1 2
timestamp 1756547599
<< locali >>
rect 635 12137 14085 12171
rect 635 11061 669 12137
rect 14051 11061 14085 12137
rect 635 11027 14085 11061
<< viali >>
rect 599 12275 14121 12309
rect 499 10989 533 12209
rect 14187 10989 14221 12209
rect 599 10889 14121 10923
<< metal1 >>
rect 878 12315 884 12318
rect 493 12309 884 12315
rect 936 12315 942 12318
rect 1394 12315 1400 12318
rect 936 12309 1400 12315
rect 1452 12315 1458 12318
rect 1910 12315 1916 12318
rect 1452 12309 1916 12315
rect 1968 12315 1974 12318
rect 2426 12315 2432 12318
rect 1968 12309 2432 12315
rect 2484 12315 2490 12318
rect 2942 12315 2948 12318
rect 2484 12309 2948 12315
rect 3000 12315 3006 12318
rect 3458 12315 3464 12318
rect 3000 12309 3464 12315
rect 3516 12315 3522 12318
rect 3974 12315 3980 12318
rect 3516 12309 3980 12315
rect 4032 12315 4038 12318
rect 4490 12315 4496 12318
rect 4032 12309 4496 12315
rect 4548 12315 4554 12318
rect 5006 12315 5012 12318
rect 4548 12309 5012 12315
rect 5064 12315 5070 12318
rect 5522 12315 5528 12318
rect 5064 12309 5528 12315
rect 5580 12315 5586 12318
rect 6038 12315 6044 12318
rect 5580 12309 6044 12315
rect 6096 12315 6102 12318
rect 6554 12315 6560 12318
rect 6096 12309 6560 12315
rect 6612 12315 6618 12318
rect 7070 12315 7076 12318
rect 6612 12309 7076 12315
rect 7128 12315 7134 12318
rect 7586 12315 7592 12318
rect 7128 12309 7592 12315
rect 7644 12315 7650 12318
rect 8102 12315 8108 12318
rect 7644 12309 8108 12315
rect 8160 12315 8166 12318
rect 8618 12315 8624 12318
rect 8160 12309 8624 12315
rect 8676 12315 8682 12318
rect 9134 12315 9140 12318
rect 8676 12309 9140 12315
rect 9192 12315 9198 12318
rect 9650 12315 9656 12318
rect 9192 12309 9656 12315
rect 9708 12315 9714 12318
rect 10166 12315 10172 12318
rect 9708 12309 10172 12315
rect 10224 12315 10230 12318
rect 10682 12315 10688 12318
rect 10224 12309 10688 12315
rect 10740 12315 10746 12318
rect 11198 12315 11204 12318
rect 10740 12309 11204 12315
rect 11256 12315 11262 12318
rect 11714 12315 11720 12318
rect 11256 12309 11720 12315
rect 11772 12315 11778 12318
rect 12230 12315 12236 12318
rect 11772 12309 12236 12315
rect 12288 12315 12294 12318
rect 12746 12315 12752 12318
rect 12288 12309 12752 12315
rect 12804 12315 12810 12318
rect 13262 12315 13268 12318
rect 12804 12309 13268 12315
rect 13320 12315 13326 12318
rect 13778 12315 13784 12318
rect 13320 12309 13784 12315
rect 13836 12315 13842 12318
rect 13836 12309 14227 12315
rect 493 12275 599 12309
rect 14121 12275 14227 12309
rect 493 12269 884 12275
rect 493 12209 539 12269
rect 878 12266 884 12269
rect 936 12269 1400 12275
rect 936 12266 942 12269
rect 1394 12266 1400 12269
rect 1452 12269 1916 12275
rect 1452 12266 1458 12269
rect 1910 12266 1916 12269
rect 1968 12269 2432 12275
rect 1968 12266 1974 12269
rect 2426 12266 2432 12269
rect 2484 12269 2948 12275
rect 2484 12266 2490 12269
rect 2942 12266 2948 12269
rect 3000 12269 3464 12275
rect 3000 12266 3006 12269
rect 3458 12266 3464 12269
rect 3516 12269 3980 12275
rect 3516 12266 3522 12269
rect 3974 12266 3980 12269
rect 4032 12269 4496 12275
rect 4032 12266 4038 12269
rect 4490 12266 4496 12269
rect 4548 12269 5012 12275
rect 4548 12266 4554 12269
rect 5006 12266 5012 12269
rect 5064 12269 5528 12275
rect 5064 12266 5070 12269
rect 5522 12266 5528 12269
rect 5580 12269 6044 12275
rect 5580 12266 5586 12269
rect 6038 12266 6044 12269
rect 6096 12269 6560 12275
rect 6096 12266 6102 12269
rect 6554 12266 6560 12269
rect 6612 12269 7076 12275
rect 6612 12266 6618 12269
rect 7070 12266 7076 12269
rect 7128 12269 7592 12275
rect 7128 12266 7134 12269
rect 7586 12266 7592 12269
rect 7644 12269 8108 12275
rect 7644 12266 7650 12269
rect 8102 12266 8108 12269
rect 8160 12269 8624 12275
rect 8160 12266 8166 12269
rect 8618 12266 8624 12269
rect 8676 12269 9140 12275
rect 8676 12266 8682 12269
rect 9134 12266 9140 12269
rect 9192 12269 9656 12275
rect 9192 12266 9198 12269
rect 9650 12266 9656 12269
rect 9708 12269 10172 12275
rect 9708 12266 9714 12269
rect 10166 12266 10172 12269
rect 10224 12269 10688 12275
rect 10224 12266 10230 12269
rect 10682 12266 10688 12269
rect 10740 12269 11204 12275
rect 10740 12266 10746 12269
rect 11198 12266 11204 12269
rect 11256 12269 11720 12275
rect 11256 12266 11262 12269
rect 11714 12266 11720 12269
rect 11772 12269 12236 12275
rect 11772 12266 11778 12269
rect 12230 12266 12236 12269
rect 12288 12269 12752 12275
rect 12288 12266 12294 12269
rect 12746 12266 12752 12269
rect 12804 12269 13268 12275
rect 12804 12266 12810 12269
rect 13262 12266 13268 12269
rect 13320 12269 13784 12275
rect 13320 12266 13326 12269
rect 13778 12266 13784 12269
rect 13836 12269 14227 12275
rect 13836 12266 13842 12269
rect 493 10989 499 12209
rect 533 10989 539 12209
rect 14181 12209 14227 12269
rect 626 12131 14094 12177
rect 626 12093 678 12131
rect 626 11293 678 11393
rect 626 11067 678 11105
rect 884 12093 936 12099
rect 884 11099 936 11105
rect 1142 12093 1194 12099
rect 1142 11099 1194 11105
rect 1400 12093 1452 12099
rect 1400 11099 1452 11105
rect 1658 12093 1710 12099
rect 1658 11099 1710 11105
rect 1916 12093 1968 12099
rect 1916 11099 1968 11105
rect 2174 12093 2226 12099
rect 2174 11099 2226 11105
rect 2432 12093 2484 12099
rect 2432 11099 2484 11105
rect 2690 12093 2742 12099
rect 2690 11099 2742 11105
rect 2948 12093 3000 12099
rect 2948 11099 3000 11105
rect 3206 12093 3258 12099
rect 3206 11099 3258 11105
rect 3464 12093 3516 12099
rect 3464 11099 3516 11105
rect 3722 12093 3774 12099
rect 3722 11099 3774 11105
rect 3980 12093 4032 12099
rect 3980 11099 4032 11105
rect 4238 12093 4290 12099
rect 4238 11099 4290 11105
rect 4496 12093 4548 12099
rect 4496 11099 4548 11105
rect 4754 12093 4806 12099
rect 4754 11099 4806 11105
rect 5012 12093 5064 12099
rect 5012 11099 5064 11105
rect 5270 12093 5322 12099
rect 5270 11099 5322 11105
rect 5528 12093 5580 12099
rect 5528 11099 5580 11105
rect 5786 12093 5838 12099
rect 5786 11099 5838 11105
rect 6044 12093 6096 12099
rect 6044 11099 6096 11105
rect 6302 12093 6354 12099
rect 6302 11099 6354 11105
rect 6560 12093 6612 12099
rect 6560 11099 6612 11105
rect 6818 12093 6870 12099
rect 6818 11099 6870 11105
rect 7076 12093 7128 12099
rect 7076 11099 7128 11105
rect 7334 12093 7386 12099
rect 7334 11099 7386 11105
rect 7592 12093 7644 12099
rect 7592 11099 7644 11105
rect 7850 12093 7902 12099
rect 7850 11099 7902 11105
rect 8108 12093 8160 12099
rect 8108 11099 8160 11105
rect 8366 12093 8418 12099
rect 8366 11099 8418 11105
rect 8624 12093 8676 12099
rect 8624 11099 8676 11105
rect 8882 12093 8934 12099
rect 8882 11099 8934 11105
rect 9140 12093 9192 12099
rect 9140 11099 9192 11105
rect 9398 12093 9450 12099
rect 9398 11099 9450 11105
rect 9656 12093 9708 12099
rect 9656 11099 9708 11105
rect 9914 12093 9966 12099
rect 9914 11099 9966 11105
rect 10172 12093 10224 12099
rect 10172 11099 10224 11105
rect 10430 12093 10482 12099
rect 10430 11099 10482 11105
rect 10688 12093 10740 12099
rect 10688 11099 10740 11105
rect 10946 12093 10998 12099
rect 10946 11099 10998 11105
rect 11204 12093 11256 12099
rect 11204 11099 11256 11105
rect 11462 12093 11514 12099
rect 11462 11099 11514 11105
rect 11720 12093 11772 12099
rect 11720 11099 11772 11105
rect 11978 12093 12030 12099
rect 11978 11099 12030 11105
rect 12236 12093 12288 12099
rect 12236 11099 12288 11105
rect 12494 12093 12546 12099
rect 12494 11099 12546 11105
rect 12752 12093 12804 12099
rect 12752 11099 12804 11105
rect 13010 12093 13062 12099
rect 13010 11099 13062 11105
rect 13268 12093 13320 12099
rect 13268 11099 13320 11105
rect 13526 12093 13578 12099
rect 13526 11099 13578 11105
rect 13784 12093 13836 12099
rect 13784 11099 13836 11105
rect 14042 12093 14094 12131
rect 14042 11067 14094 11105
rect 626 11021 14094 11067
rect 493 10929 539 10989
rect 14181 10989 14187 12209
rect 14221 10989 14227 12209
rect 878 10929 884 10932
rect 493 10923 884 10929
rect 936 10929 942 10932
rect 1394 10929 1400 10932
rect 936 10923 1400 10929
rect 1452 10929 1458 10932
rect 1910 10929 1916 10932
rect 1452 10923 1916 10929
rect 1968 10929 1974 10932
rect 2426 10929 2432 10932
rect 1968 10923 2432 10929
rect 2484 10929 2490 10932
rect 2942 10929 2948 10932
rect 2484 10923 2948 10929
rect 3000 10929 3006 10932
rect 3458 10929 3464 10932
rect 3000 10923 3464 10929
rect 3516 10929 3522 10932
rect 3974 10929 3980 10932
rect 3516 10923 3980 10929
rect 4032 10929 4038 10932
rect 4490 10929 4496 10932
rect 4032 10923 4496 10929
rect 4548 10929 4554 10932
rect 5006 10929 5012 10932
rect 4548 10923 5012 10929
rect 5064 10929 5070 10932
rect 5522 10929 5528 10932
rect 5064 10923 5528 10929
rect 5580 10929 5586 10932
rect 6038 10929 6044 10932
rect 5580 10923 6044 10929
rect 6096 10929 6102 10932
rect 6554 10929 6560 10932
rect 6096 10923 6560 10929
rect 6612 10929 6618 10932
rect 7070 10929 7076 10932
rect 6612 10923 7076 10929
rect 7128 10929 7134 10932
rect 7586 10929 7592 10932
rect 7128 10923 7592 10929
rect 7644 10929 7650 10932
rect 8102 10929 8108 10932
rect 7644 10923 8108 10929
rect 8160 10929 8166 10932
rect 8618 10929 8624 10932
rect 8160 10923 8624 10929
rect 8676 10929 8682 10932
rect 9134 10929 9140 10932
rect 8676 10923 9140 10929
rect 9192 10929 9198 10932
rect 9650 10929 9656 10932
rect 9192 10923 9656 10929
rect 9708 10929 9714 10932
rect 10166 10929 10172 10932
rect 9708 10923 10172 10929
rect 10224 10929 10230 10932
rect 10682 10929 10688 10932
rect 10224 10923 10688 10929
rect 10740 10929 10746 10932
rect 11198 10929 11204 10932
rect 10740 10923 11204 10929
rect 11256 10929 11262 10932
rect 11714 10929 11720 10932
rect 11256 10923 11720 10929
rect 11772 10929 11778 10932
rect 12230 10929 12236 10932
rect 11772 10923 12236 10929
rect 12288 10929 12294 10932
rect 12746 10929 12752 10932
rect 12288 10923 12752 10929
rect 12804 10929 12810 10932
rect 13262 10929 13268 10932
rect 12804 10923 13268 10929
rect 13320 10929 13326 10932
rect 13778 10929 13784 10932
rect 13320 10923 13784 10929
rect 13836 10929 13842 10932
rect 14181 10929 14227 10989
rect 13836 10923 14227 10929
rect 493 10889 599 10923
rect 14121 10889 14227 10923
rect 493 10883 884 10889
rect 878 10880 884 10883
rect 936 10883 1400 10889
rect 936 10880 942 10883
rect 1394 10880 1400 10883
rect 1452 10883 1916 10889
rect 1452 10880 1458 10883
rect 1910 10880 1916 10883
rect 1968 10883 2432 10889
rect 1968 10880 1974 10883
rect 2426 10880 2432 10883
rect 2484 10883 2948 10889
rect 2484 10880 2490 10883
rect 2942 10880 2948 10883
rect 3000 10883 3464 10889
rect 3000 10880 3006 10883
rect 3458 10880 3464 10883
rect 3516 10883 3980 10889
rect 3516 10880 3522 10883
rect 3974 10880 3980 10883
rect 4032 10883 4496 10889
rect 4032 10880 4038 10883
rect 4490 10880 4496 10883
rect 4548 10883 5012 10889
rect 4548 10880 4554 10883
rect 5006 10880 5012 10883
rect 5064 10883 5528 10889
rect 5064 10880 5070 10883
rect 5522 10880 5528 10883
rect 5580 10883 6044 10889
rect 5580 10880 5586 10883
rect 6038 10880 6044 10883
rect 6096 10883 6560 10889
rect 6096 10880 6102 10883
rect 6554 10880 6560 10883
rect 6612 10883 7076 10889
rect 6612 10880 6618 10883
rect 7070 10880 7076 10883
rect 7128 10883 7592 10889
rect 7128 10880 7134 10883
rect 7586 10880 7592 10883
rect 7644 10883 8108 10889
rect 7644 10880 7650 10883
rect 8102 10880 8108 10883
rect 8160 10883 8624 10889
rect 8160 10880 8166 10883
rect 8618 10880 8624 10883
rect 8676 10883 9140 10889
rect 8676 10880 8682 10883
rect 9134 10880 9140 10883
rect 9192 10883 9656 10889
rect 9192 10880 9198 10883
rect 9650 10880 9656 10883
rect 9708 10883 10172 10889
rect 9708 10880 9714 10883
rect 10166 10880 10172 10883
rect 10224 10883 10688 10889
rect 10224 10880 10230 10883
rect 10682 10880 10688 10883
rect 10740 10883 11204 10889
rect 10740 10880 10746 10883
rect 11198 10880 11204 10883
rect 11256 10883 11720 10889
rect 11256 10880 11262 10883
rect 11714 10880 11720 10883
rect 11772 10883 12236 10889
rect 11772 10880 11778 10883
rect 12230 10880 12236 10883
rect 12288 10883 12752 10889
rect 12288 10880 12294 10883
rect 12746 10880 12752 10883
rect 12804 10883 13268 10889
rect 12804 10880 12810 10883
rect 13262 10880 13268 10883
rect 13320 10883 13784 10889
rect 13320 10880 13326 10883
rect 13778 10880 13784 10883
rect 13836 10883 14227 10889
rect 13836 10880 13842 10883
<< via1 >>
rect 884 12309 936 12318
rect 1400 12309 1452 12318
rect 1916 12309 1968 12318
rect 2432 12309 2484 12318
rect 2948 12309 3000 12318
rect 3464 12309 3516 12318
rect 3980 12309 4032 12318
rect 4496 12309 4548 12318
rect 5012 12309 5064 12318
rect 5528 12309 5580 12318
rect 6044 12309 6096 12318
rect 6560 12309 6612 12318
rect 7076 12309 7128 12318
rect 7592 12309 7644 12318
rect 8108 12309 8160 12318
rect 8624 12309 8676 12318
rect 9140 12309 9192 12318
rect 9656 12309 9708 12318
rect 10172 12309 10224 12318
rect 10688 12309 10740 12318
rect 11204 12309 11256 12318
rect 11720 12309 11772 12318
rect 12236 12309 12288 12318
rect 12752 12309 12804 12318
rect 13268 12309 13320 12318
rect 13784 12309 13836 12318
rect 884 12275 936 12309
rect 1400 12275 1452 12309
rect 1916 12275 1968 12309
rect 2432 12275 2484 12309
rect 2948 12275 3000 12309
rect 3464 12275 3516 12309
rect 3980 12275 4032 12309
rect 4496 12275 4548 12309
rect 5012 12275 5064 12309
rect 5528 12275 5580 12309
rect 6044 12275 6096 12309
rect 6560 12275 6612 12309
rect 7076 12275 7128 12309
rect 7592 12275 7644 12309
rect 8108 12275 8160 12309
rect 8624 12275 8676 12309
rect 9140 12275 9192 12309
rect 9656 12275 9708 12309
rect 10172 12275 10224 12309
rect 10688 12275 10740 12309
rect 11204 12275 11256 12309
rect 11720 12275 11772 12309
rect 12236 12275 12288 12309
rect 12752 12275 12804 12309
rect 13268 12275 13320 12309
rect 13784 12275 13836 12309
rect 884 12266 936 12275
rect 1400 12266 1452 12275
rect 1916 12266 1968 12275
rect 2432 12266 2484 12275
rect 2948 12266 3000 12275
rect 3464 12266 3516 12275
rect 3980 12266 4032 12275
rect 4496 12266 4548 12275
rect 5012 12266 5064 12275
rect 5528 12266 5580 12275
rect 6044 12266 6096 12275
rect 6560 12266 6612 12275
rect 7076 12266 7128 12275
rect 7592 12266 7644 12275
rect 8108 12266 8160 12275
rect 8624 12266 8676 12275
rect 9140 12266 9192 12275
rect 9656 12266 9708 12275
rect 10172 12266 10224 12275
rect 10688 12266 10740 12275
rect 11204 12266 11256 12275
rect 11720 12266 11772 12275
rect 12236 12266 12288 12275
rect 12752 12266 12804 12275
rect 13268 12266 13320 12275
rect 13784 12266 13836 12275
rect 626 11393 678 12093
rect 626 11105 678 11293
rect 884 11105 936 12093
rect 1142 11105 1194 12093
rect 1400 11105 1452 12093
rect 1658 11105 1710 12093
rect 1916 11105 1968 12093
rect 2174 11105 2226 12093
rect 2432 11105 2484 12093
rect 2690 11105 2742 12093
rect 2948 11105 3000 12093
rect 3206 11105 3258 12093
rect 3464 11105 3516 12093
rect 3722 11105 3774 12093
rect 3980 11105 4032 12093
rect 4238 11105 4290 12093
rect 4496 11105 4548 12093
rect 4754 11105 4806 12093
rect 5012 11105 5064 12093
rect 5270 11105 5322 12093
rect 5528 11105 5580 12093
rect 5786 11105 5838 12093
rect 6044 11105 6096 12093
rect 6302 11105 6354 12093
rect 6560 11105 6612 12093
rect 6818 11105 6870 12093
rect 7076 11105 7128 12093
rect 7334 11105 7386 12093
rect 7592 11105 7644 12093
rect 7850 11105 7902 12093
rect 8108 11105 8160 12093
rect 8366 11105 8418 12093
rect 8624 11105 8676 12093
rect 8882 11105 8934 12093
rect 9140 11105 9192 12093
rect 9398 11105 9450 12093
rect 9656 11105 9708 12093
rect 9914 11105 9966 12093
rect 10172 11105 10224 12093
rect 10430 11105 10482 12093
rect 10688 11105 10740 12093
rect 10946 11105 10998 12093
rect 11204 11105 11256 12093
rect 11462 11105 11514 12093
rect 11720 11105 11772 12093
rect 11978 11105 12030 12093
rect 12236 11105 12288 12093
rect 12494 11105 12546 12093
rect 12752 11105 12804 12093
rect 13010 11105 13062 12093
rect 13268 11105 13320 12093
rect 13526 11105 13578 12093
rect 13784 11105 13836 12093
rect 14042 11105 14094 12093
rect 884 10923 936 10932
rect 1400 10923 1452 10932
rect 1916 10923 1968 10932
rect 2432 10923 2484 10932
rect 2948 10923 3000 10932
rect 3464 10923 3516 10932
rect 3980 10923 4032 10932
rect 4496 10923 4548 10932
rect 5012 10923 5064 10932
rect 5528 10923 5580 10932
rect 6044 10923 6096 10932
rect 6560 10923 6612 10932
rect 7076 10923 7128 10932
rect 7592 10923 7644 10932
rect 8108 10923 8160 10932
rect 8624 10923 8676 10932
rect 9140 10923 9192 10932
rect 9656 10923 9708 10932
rect 10172 10923 10224 10932
rect 10688 10923 10740 10932
rect 11204 10923 11256 10932
rect 11720 10923 11772 10932
rect 12236 10923 12288 10932
rect 12752 10923 12804 10932
rect 13268 10923 13320 10932
rect 13784 10923 13836 10932
rect 884 10889 936 10923
rect 1400 10889 1452 10923
rect 1916 10889 1968 10923
rect 2432 10889 2484 10923
rect 2948 10889 3000 10923
rect 3464 10889 3516 10923
rect 3980 10889 4032 10923
rect 4496 10889 4548 10923
rect 5012 10889 5064 10923
rect 5528 10889 5580 10923
rect 6044 10889 6096 10923
rect 6560 10889 6612 10923
rect 7076 10889 7128 10923
rect 7592 10889 7644 10923
rect 8108 10889 8160 10923
rect 8624 10889 8676 10923
rect 9140 10889 9192 10923
rect 9656 10889 9708 10923
rect 10172 10889 10224 10923
rect 10688 10889 10740 10923
rect 11204 10889 11256 10923
rect 11720 10889 11772 10923
rect 12236 10889 12288 10923
rect 12752 10889 12804 10923
rect 13268 10889 13320 10923
rect 13784 10889 13836 10923
rect 884 10880 936 10889
rect 1400 10880 1452 10889
rect 1916 10880 1968 10889
rect 2432 10880 2484 10889
rect 2948 10880 3000 10889
rect 3464 10880 3516 10889
rect 3980 10880 4032 10889
rect 4496 10880 4548 10889
rect 5012 10880 5064 10889
rect 5528 10880 5580 10889
rect 6044 10880 6096 10889
rect 6560 10880 6612 10889
rect 7076 10880 7128 10889
rect 7592 10880 7644 10889
rect 8108 10880 8160 10889
rect 8624 10880 8676 10889
rect 9140 10880 9192 10889
rect 9656 10880 9708 10889
rect 10172 10880 10224 10889
rect 10688 10880 10740 10889
rect 11204 10880 11256 10889
rect 11720 10880 11772 10889
rect 12236 10880 12288 10889
rect 12752 10880 12804 10889
rect 13268 10880 13320 10889
rect 13784 10880 13836 10889
<< metal2 >>
rect 626 12093 678 12923
rect 1142 12753 1194 12923
rect 1060 12744 1276 12753
rect 1060 12653 1276 12662
rect 878 12266 884 12318
rect 936 12266 942 12318
rect 884 12093 936 12266
rect 842 11728 884 11737
rect 1142 12093 1194 12653
rect 1658 12583 1710 12923
rect 1576 12574 1792 12583
rect 1576 12483 1792 12492
rect 1394 12266 1400 12318
rect 1452 12266 1458 12318
rect 936 11728 978 11737
rect 842 11459 884 11468
rect 626 11293 678 11393
rect 626 10373 678 11105
rect 936 11459 978 11468
rect 884 10932 936 11105
rect 1400 12093 1452 12266
rect 1358 11728 1400 11737
rect 1658 12093 1710 12483
rect 1910 12266 1916 12318
rect 1968 12266 1974 12318
rect 1452 11728 1494 11737
rect 1358 11459 1400 11468
rect 878 10880 884 10932
rect 936 10880 942 10932
rect 544 10364 760 10373
rect 544 10273 760 10282
rect 1142 10273 1194 11105
rect 1452 11459 1494 11468
rect 1400 10932 1452 11105
rect 1916 12093 1968 12266
rect 2174 12243 2226 12923
rect 2426 12266 2432 12318
rect 2484 12266 2490 12318
rect 2092 12234 2308 12243
rect 2092 12143 2308 12152
rect 1874 11728 1916 11737
rect 2174 12093 2226 12143
rect 1968 11728 2010 11737
rect 1874 11459 1916 11468
rect 1394 10880 1400 10932
rect 1452 10880 1458 10932
rect 1658 10273 1710 11105
rect 1968 11459 2010 11468
rect 1916 10932 1968 11105
rect 2432 12093 2484 12266
rect 2390 11728 2432 11737
rect 2690 12093 2742 12923
rect 3206 12413 3258 12923
rect 3124 12404 3340 12413
rect 2942 12266 2948 12318
rect 3000 12266 3006 12318
rect 3124 12313 3340 12322
rect 2484 11728 2526 11737
rect 2390 11459 2432 11468
rect 1910 10880 1916 10932
rect 1968 10880 1974 10932
rect 2174 10273 2226 11105
rect 2484 11459 2526 11468
rect 2432 10932 2484 11105
rect 2948 12093 3000 12266
rect 2906 11728 2948 11737
rect 3206 12093 3258 12313
rect 3458 12266 3464 12318
rect 3516 12266 3522 12318
rect 3000 11728 3042 11737
rect 2906 11459 2948 11468
rect 2426 10880 2432 10932
rect 2484 10880 2490 10932
rect 2690 10883 2742 11105
rect 3000 11459 3042 11468
rect 2948 10932 3000 11105
rect 3464 12093 3516 12266
rect 3422 11728 3464 11737
rect 3722 12093 3774 12923
rect 3974 12266 3980 12318
rect 4032 12266 4038 12318
rect 3640 12064 3722 12073
rect 3980 12093 4032 12266
rect 3774 12064 3856 12073
rect 3640 11973 3722 11982
rect 3516 11728 3558 11737
rect 3422 11459 3464 11468
rect 2608 10874 2824 10883
rect 2942 10880 2948 10932
rect 3000 10880 3006 10932
rect 2608 10783 2824 10792
rect 2690 10273 2742 10783
rect 3206 10273 3258 11105
rect 3516 11459 3558 11468
rect 3464 10932 3516 11105
rect 3774 11973 3856 11982
rect 3938 11728 3980 11737
rect 4238 12093 4290 12923
rect 4490 12266 4496 12318
rect 4548 12266 4554 12318
rect 4156 12064 4238 12073
rect 4496 12093 4548 12266
rect 4290 12064 4372 12073
rect 4156 11973 4238 11982
rect 4032 11728 4074 11737
rect 3938 11459 3980 11468
rect 3458 10880 3464 10932
rect 3516 10880 3522 10932
rect 3722 10273 3774 11105
rect 4032 11459 4074 11468
rect 3980 10932 4032 11105
rect 4290 11973 4372 11982
rect 4454 11728 4496 11737
rect 4754 12093 4806 12923
rect 5006 12266 5012 12318
rect 5064 12266 5070 12318
rect 4548 11728 4590 11737
rect 4454 11459 4496 11468
rect 3974 10880 3980 10932
rect 4032 10880 4038 10932
rect 4238 10273 4290 11105
rect 4548 11459 4590 11468
rect 4672 11214 4754 11223
rect 5012 12093 5064 12266
rect 4970 11728 5012 11737
rect 5270 12093 5322 12923
rect 5522 12266 5528 12318
rect 5580 12266 5586 12318
rect 5064 11728 5106 11737
rect 4970 11459 5012 11468
rect 4806 11214 4888 11223
rect 4672 11123 4754 11132
rect 4496 10932 4548 11105
rect 4806 11123 4888 11132
rect 4490 10880 4496 10932
rect 4548 10880 4554 10932
rect 4754 10273 4806 11105
rect 5064 11459 5106 11468
rect 5188 11214 5270 11223
rect 5528 12093 5580 12266
rect 5486 11728 5528 11737
rect 5786 12093 5838 12923
rect 6038 12266 6044 12318
rect 6096 12266 6102 12318
rect 5580 11728 5622 11737
rect 5486 11459 5528 11468
rect 5322 11214 5404 11223
rect 5188 11123 5270 11132
rect 5012 10932 5064 11105
rect 5322 11123 5404 11132
rect 5006 10880 5012 10932
rect 5064 10880 5070 10932
rect 5270 10273 5322 11105
rect 5580 11459 5622 11468
rect 5528 10932 5580 11105
rect 6044 12093 6096 12266
rect 6002 11728 6044 11737
rect 6302 12093 6354 12923
rect 6554 12266 6560 12318
rect 6612 12266 6618 12318
rect 6096 11728 6138 11737
rect 6002 11459 6044 11468
rect 5786 11053 5838 11105
rect 6096 11459 6138 11468
rect 6220 11384 6302 11393
rect 6560 12093 6612 12266
rect 6518 11728 6560 11737
rect 6818 12093 6870 12923
rect 7252 12914 7468 12923
rect 7252 12823 7468 12832
rect 7070 12266 7076 12318
rect 7128 12266 7134 12318
rect 6736 11894 6818 11903
rect 7076 12093 7128 12266
rect 6870 11894 6952 11903
rect 6736 11803 6818 11812
rect 6612 11728 6654 11737
rect 6518 11459 6560 11468
rect 6354 11384 6436 11393
rect 6220 11293 6302 11302
rect 5704 11044 5920 11053
rect 5704 10953 5920 10962
rect 5522 10880 5528 10932
rect 5580 10880 5586 10932
rect 5786 10273 5838 10953
rect 6044 10932 6096 11105
rect 6354 11293 6436 11302
rect 6038 10880 6044 10932
rect 6096 10880 6102 10932
rect 6302 10273 6354 11105
rect 6612 11459 6654 11468
rect 6560 10932 6612 11105
rect 6870 11803 6952 11812
rect 7034 11728 7076 11737
rect 7334 12093 7386 12823
rect 7586 12266 7592 12318
rect 7644 12266 7650 12318
rect 7128 11728 7170 11737
rect 7034 11459 7076 11468
rect 6554 10880 6560 10932
rect 6612 10880 6618 10932
rect 6818 10273 6870 11105
rect 7128 11459 7170 11468
rect 7076 10932 7128 11105
rect 7592 12093 7644 12266
rect 7550 11728 7592 11737
rect 7850 12093 7902 12923
rect 8102 12266 8108 12318
rect 8160 12266 8166 12318
rect 7768 11894 7850 11903
rect 8108 12093 8160 12266
rect 7902 11894 7984 11903
rect 7768 11803 7850 11812
rect 7644 11728 7686 11737
rect 7550 11459 7592 11468
rect 7070 10880 7076 10932
rect 7128 10880 7134 10932
rect 7334 10273 7386 11105
rect 7644 11459 7686 11468
rect 7592 10932 7644 11105
rect 7902 11803 7984 11812
rect 8066 11728 8108 11737
rect 8366 12093 8418 12923
rect 8618 12266 8624 12318
rect 8676 12266 8682 12318
rect 8160 11728 8202 11737
rect 8066 11459 8108 11468
rect 7586 10880 7592 10932
rect 7644 10880 7650 10932
rect 7850 10273 7902 11105
rect 8160 11459 8202 11468
rect 8284 11384 8366 11393
rect 8624 12093 8676 12266
rect 8582 11728 8624 11737
rect 8882 12093 8934 12923
rect 9134 12266 9140 12318
rect 9192 12266 9198 12318
rect 8676 11728 8718 11737
rect 8582 11459 8624 11468
rect 8418 11384 8500 11393
rect 8284 11293 8366 11302
rect 8108 10932 8160 11105
rect 8418 11293 8500 11302
rect 8102 10880 8108 10932
rect 8160 10880 8166 10932
rect 8366 10273 8418 11105
rect 8676 11459 8718 11468
rect 8624 10932 8676 11105
rect 9140 12093 9192 12266
rect 9098 11728 9140 11737
rect 9398 12093 9450 12923
rect 9650 12266 9656 12318
rect 9708 12266 9714 12318
rect 9192 11728 9234 11737
rect 9098 11459 9140 11468
rect 8882 11053 8934 11105
rect 9192 11459 9234 11468
rect 9316 11214 9398 11223
rect 9656 12093 9708 12266
rect 9614 11728 9656 11737
rect 9914 12093 9966 12923
rect 10166 12266 10172 12318
rect 10224 12266 10230 12318
rect 9708 11728 9750 11737
rect 9614 11459 9656 11468
rect 9450 11214 9532 11223
rect 9316 11123 9398 11132
rect 8800 11044 9016 11053
rect 8800 10953 9016 10962
rect 8618 10880 8624 10932
rect 8676 10880 8682 10932
rect 8882 10273 8934 10953
rect 9140 10932 9192 11105
rect 9450 11123 9532 11132
rect 9134 10880 9140 10932
rect 9192 10880 9198 10932
rect 9398 10273 9450 11105
rect 9708 11459 9750 11468
rect 9832 11214 9914 11223
rect 10172 12093 10224 12266
rect 10130 11728 10172 11737
rect 10430 12093 10482 12923
rect 10682 12266 10688 12318
rect 10740 12266 10746 12318
rect 10348 12064 10430 12073
rect 10688 12093 10740 12266
rect 10482 12064 10564 12073
rect 10348 11973 10430 11982
rect 10224 11728 10266 11737
rect 10130 11459 10172 11468
rect 9966 11214 10048 11223
rect 9832 11123 9914 11132
rect 9656 10932 9708 11105
rect 9966 11123 10048 11132
rect 9650 10880 9656 10932
rect 9708 10880 9714 10932
rect 9914 10273 9966 11105
rect 10224 11459 10266 11468
rect 10172 10932 10224 11105
rect 10482 11973 10564 11982
rect 10646 11728 10688 11737
rect 10946 12093 10998 12923
rect 11462 12413 11514 12923
rect 11380 12404 11596 12413
rect 11198 12266 11204 12318
rect 11256 12266 11262 12318
rect 11380 12313 11596 12322
rect 10864 12064 10946 12073
rect 11204 12093 11256 12266
rect 10998 12064 11080 12073
rect 10864 11973 10946 11982
rect 10740 11728 10782 11737
rect 10646 11459 10688 11468
rect 10166 10880 10172 10932
rect 10224 10880 10230 10932
rect 10430 10273 10482 11105
rect 10740 11459 10782 11468
rect 10688 10932 10740 11105
rect 10998 11973 11080 11982
rect 11162 11728 11204 11737
rect 11462 12093 11514 12313
rect 11714 12266 11720 12318
rect 11772 12266 11778 12318
rect 11256 11728 11298 11737
rect 11162 11459 11204 11468
rect 10682 10880 10688 10932
rect 10740 10880 10746 10932
rect 10946 10273 10998 11105
rect 11256 11459 11298 11468
rect 11204 10932 11256 11105
rect 11720 12093 11772 12266
rect 11678 11728 11720 11737
rect 11978 12093 12030 12923
rect 12230 12266 12236 12318
rect 12288 12266 12294 12318
rect 11772 11728 11814 11737
rect 11678 11459 11720 11468
rect 11198 10880 11204 10932
rect 11256 10880 11262 10932
rect 11462 10273 11514 11105
rect 11772 11459 11814 11468
rect 11720 10932 11772 11105
rect 12236 12093 12288 12266
rect 12494 12243 12546 12923
rect 12746 12266 12752 12318
rect 12804 12266 12810 12318
rect 12412 12234 12628 12243
rect 12412 12143 12628 12152
rect 12194 11728 12236 11737
rect 12494 12093 12546 12143
rect 12288 11728 12330 11737
rect 12194 11459 12236 11468
rect 11714 10880 11720 10932
rect 11772 10880 11778 10932
rect 11978 10883 12030 11105
rect 12288 11459 12330 11468
rect 12236 10932 12288 11105
rect 12752 12093 12804 12266
rect 12710 11728 12752 11737
rect 13010 12093 13062 12923
rect 13262 12266 13268 12318
rect 13320 12266 13326 12318
rect 12804 11728 12846 11737
rect 12710 11459 12752 11468
rect 11896 10874 12112 10883
rect 12230 10880 12236 10932
rect 12288 10880 12294 10932
rect 11896 10783 12112 10792
rect 11978 10273 12030 10783
rect 12494 10273 12546 11105
rect 12804 11459 12846 11468
rect 12752 10932 12804 11105
rect 13268 12093 13320 12266
rect 13226 11728 13268 11737
rect 13526 12093 13578 12923
rect 13778 12266 13784 12318
rect 13836 12266 13842 12318
rect 13320 11728 13362 11737
rect 13226 11459 13268 11468
rect 12746 10880 12752 10932
rect 12804 10880 12810 10932
rect 13010 10713 13062 11105
rect 13320 11459 13362 11468
rect 13268 10932 13320 11105
rect 13784 12093 13836 12266
rect 13742 11728 13784 11737
rect 14042 12093 14094 12923
rect 13836 11728 13878 11737
rect 13742 11459 13784 11468
rect 13262 10880 13268 10932
rect 13320 10880 13326 10932
rect 12928 10704 13144 10713
rect 12928 10613 13144 10622
rect 13010 10273 13062 10613
rect 13526 10543 13578 11105
rect 13836 11459 13878 11468
rect 13784 10932 13836 11105
rect 13778 10880 13784 10932
rect 13836 10880 13842 10932
rect 13444 10534 13660 10543
rect 13444 10443 13660 10452
rect 13526 10273 13578 10443
rect 14042 10373 14094 11105
rect 13960 10364 14176 10373
rect 13960 10273 14176 10282
<< via2 >>
rect 1060 12662 1276 12744
rect 1576 12492 1792 12574
rect 842 11468 884 11728
rect 884 11468 936 11728
rect 936 11468 978 11728
rect 1358 11468 1400 11728
rect 1400 11468 1452 11728
rect 1452 11468 1494 11728
rect 544 10282 760 10364
rect 2092 12152 2308 12234
rect 1874 11468 1916 11728
rect 1916 11468 1968 11728
rect 1968 11468 2010 11728
rect 3124 12322 3340 12404
rect 2390 11468 2432 11728
rect 2432 11468 2484 11728
rect 2484 11468 2526 11728
rect 2906 11468 2948 11728
rect 2948 11468 3000 11728
rect 3000 11468 3042 11728
rect 3640 11982 3722 12064
rect 3722 11982 3774 12064
rect 3774 11982 3856 12064
rect 3422 11468 3464 11728
rect 3464 11468 3516 11728
rect 3516 11468 3558 11728
rect 2608 10792 2824 10874
rect 4156 11982 4238 12064
rect 4238 11982 4290 12064
rect 4290 11982 4372 12064
rect 3938 11468 3980 11728
rect 3980 11468 4032 11728
rect 4032 11468 4074 11728
rect 4454 11468 4496 11728
rect 4496 11468 4548 11728
rect 4548 11468 4590 11728
rect 4970 11468 5012 11728
rect 5012 11468 5064 11728
rect 5064 11468 5106 11728
rect 4672 11132 4754 11214
rect 4754 11132 4806 11214
rect 4806 11132 4888 11214
rect 5486 11468 5528 11728
rect 5528 11468 5580 11728
rect 5580 11468 5622 11728
rect 5188 11132 5270 11214
rect 5270 11132 5322 11214
rect 5322 11132 5404 11214
rect 6002 11468 6044 11728
rect 6044 11468 6096 11728
rect 6096 11468 6138 11728
rect 7252 12832 7468 12914
rect 6736 11812 6818 11894
rect 6818 11812 6870 11894
rect 6870 11812 6952 11894
rect 6518 11468 6560 11728
rect 6560 11468 6612 11728
rect 6612 11468 6654 11728
rect 6220 11302 6302 11384
rect 6302 11302 6354 11384
rect 6354 11302 6436 11384
rect 5704 10962 5920 11044
rect 7034 11468 7076 11728
rect 7076 11468 7128 11728
rect 7128 11468 7170 11728
rect 7768 11812 7850 11894
rect 7850 11812 7902 11894
rect 7902 11812 7984 11894
rect 7550 11468 7592 11728
rect 7592 11468 7644 11728
rect 7644 11468 7686 11728
rect 8066 11468 8108 11728
rect 8108 11468 8160 11728
rect 8160 11468 8202 11728
rect 8582 11468 8624 11728
rect 8624 11468 8676 11728
rect 8676 11468 8718 11728
rect 8284 11302 8366 11384
rect 8366 11302 8418 11384
rect 8418 11302 8500 11384
rect 9098 11468 9140 11728
rect 9140 11468 9192 11728
rect 9192 11468 9234 11728
rect 9614 11468 9656 11728
rect 9656 11468 9708 11728
rect 9708 11468 9750 11728
rect 9316 11132 9398 11214
rect 9398 11132 9450 11214
rect 9450 11132 9532 11214
rect 8800 10962 9016 11044
rect 10348 11982 10430 12064
rect 10430 11982 10482 12064
rect 10482 11982 10564 12064
rect 10130 11468 10172 11728
rect 10172 11468 10224 11728
rect 10224 11468 10266 11728
rect 9832 11132 9914 11214
rect 9914 11132 9966 11214
rect 9966 11132 10048 11214
rect 11380 12322 11596 12404
rect 10864 11982 10946 12064
rect 10946 11982 10998 12064
rect 10998 11982 11080 12064
rect 10646 11468 10688 11728
rect 10688 11468 10740 11728
rect 10740 11468 10782 11728
rect 11162 11468 11204 11728
rect 11204 11468 11256 11728
rect 11256 11468 11298 11728
rect 11678 11468 11720 11728
rect 11720 11468 11772 11728
rect 11772 11468 11814 11728
rect 12412 12152 12628 12234
rect 12194 11468 12236 11728
rect 12236 11468 12288 11728
rect 12288 11468 12330 11728
rect 12710 11468 12752 11728
rect 12752 11468 12804 11728
rect 12804 11468 12846 11728
rect 11896 10792 12112 10874
rect 13226 11468 13268 11728
rect 13268 11468 13320 11728
rect 13320 11468 13362 11728
rect 13742 11468 13784 11728
rect 13784 11468 13836 11728
rect 13836 11468 13878 11728
rect 12928 10622 13144 10704
rect 13444 10452 13660 10534
rect 13960 10282 14176 10364
<< metal3 >>
rect 20 12914 14500 12923
rect 20 12832 7252 12914
rect 7468 12832 14500 12914
rect 20 12823 14500 12832
rect 20 12752 14500 12753
rect 20 12744 9051 12752
rect 20 12662 1060 12744
rect 1276 12662 9051 12744
rect 20 12654 9051 12662
rect 9349 12654 14500 12752
rect 20 12653 14500 12654
rect 20 12582 14500 12583
rect 20 12574 13931 12582
rect 20 12492 1576 12574
rect 1792 12492 13931 12574
rect 20 12484 13931 12492
rect 14229 12484 14500 12582
rect 20 12483 14500 12484
rect 20 12412 14500 12413
rect 20 12404 6571 12412
rect 20 12322 3124 12404
rect 3340 12322 6571 12404
rect 20 12314 6571 12322
rect 6869 12404 14500 12412
rect 6869 12322 11380 12404
rect 11596 12322 14500 12404
rect 6869 12314 14500 12322
rect 20 12313 14500 12314
rect 20 12242 14500 12243
rect 20 12144 1691 12242
rect 1989 12234 14500 12242
rect 1989 12152 2092 12234
rect 2308 12152 12412 12234
rect 12628 12152 14500 12234
rect 1989 12144 14500 12152
rect 20 12143 14500 12144
rect 20 12072 14500 12073
rect 20 11974 2291 12072
rect 2589 12064 14500 12072
rect 2589 11982 3640 12064
rect 3856 11982 4156 12064
rect 4372 11982 10348 12064
rect 10564 11982 10864 12064
rect 11080 11982 14500 12064
rect 2589 11974 14500 11982
rect 20 11973 14500 11974
rect 20 11902 14500 11903
rect 20 11894 9651 11902
rect 20 11812 6736 11894
rect 6952 11812 7768 11894
rect 7984 11812 9651 11894
rect 20 11804 9651 11812
rect 9949 11804 14500 11902
rect 20 11803 14500 11804
rect 20 11732 14500 11733
rect 20 11464 341 11732
rect 579 11728 4021 11732
rect 4259 11728 7701 11732
rect 579 11468 842 11728
rect 978 11468 1358 11728
rect 1494 11468 1874 11728
rect 2010 11468 2390 11728
rect 2526 11468 2906 11728
rect 3042 11468 3422 11728
rect 3558 11468 3938 11728
rect 4259 11468 4454 11728
rect 4590 11468 4970 11728
rect 5106 11468 5486 11728
rect 5622 11468 6002 11728
rect 6138 11468 6518 11728
rect 6654 11468 7034 11728
rect 7170 11468 7550 11728
rect 7686 11468 7701 11728
rect 579 11464 4021 11468
rect 4259 11464 7701 11468
rect 7939 11728 11381 11732
rect 7939 11468 8066 11728
rect 8202 11468 8582 11728
rect 8718 11468 9098 11728
rect 9234 11468 9614 11728
rect 9750 11468 10130 11728
rect 10266 11468 10646 11728
rect 10782 11468 11162 11728
rect 11298 11468 11381 11728
rect 7939 11464 11381 11468
rect 11619 11728 14500 11732
rect 11619 11468 11678 11728
rect 11814 11468 12194 11728
rect 12330 11468 12710 11728
rect 12846 11468 13226 11728
rect 13362 11468 13742 11728
rect 13878 11468 14500 11728
rect 11619 11464 14500 11468
rect 20 11463 14500 11464
rect 20 11392 14500 11393
rect 20 11384 13331 11392
rect 20 11302 6220 11384
rect 6436 11302 8284 11384
rect 8500 11302 13331 11384
rect 20 11294 13331 11302
rect 13629 11294 14500 11392
rect 20 11293 14500 11294
rect 20 11222 14500 11223
rect 20 11214 5971 11222
rect 20 11132 4672 11214
rect 4888 11132 5188 11214
rect 5404 11132 5971 11214
rect 20 11124 5971 11132
rect 6269 11214 14500 11222
rect 6269 11132 9316 11214
rect 9532 11132 9832 11214
rect 10048 11132 14500 11214
rect 6269 11124 14500 11132
rect 20 11123 14500 11124
rect 20 11052 14500 11053
rect 20 10954 2891 11052
rect 3189 11044 14500 11052
rect 3189 10962 5704 11044
rect 5920 10962 8800 11044
rect 9016 10962 14500 11044
rect 3189 10954 14500 10962
rect 20 10953 14500 10954
rect 20 10882 14500 10883
rect 20 10874 5371 10882
rect 20 10792 2608 10874
rect 2824 10792 5371 10874
rect 20 10784 5371 10792
rect 5669 10874 14500 10882
rect 5669 10792 11896 10874
rect 12112 10792 14500 10874
rect 5669 10784 14500 10792
rect 20 10783 14500 10784
rect 20 10712 14500 10713
rect 20 10614 12731 10712
rect 13029 10704 14500 10712
rect 13144 10622 14500 10704
rect 13029 10614 14500 10622
rect 20 10613 14500 10614
rect 20 10542 14500 10543
rect 20 10444 10251 10542
rect 10549 10534 14500 10542
rect 10549 10452 13444 10534
rect 13660 10452 14500 10534
rect 10549 10444 14500 10452
rect 20 10443 14500 10444
rect 20 10364 14500 10373
rect 20 10282 544 10364
rect 760 10282 13960 10364
rect 14176 10282 14500 10364
rect 20 10273 14500 10282
rect 954 5846 1001 5910
rect 1065 5846 1071 5910
rect 4634 5846 4681 5910
rect 4745 5846 4751 5910
rect 8314 5846 8361 5910
rect 8425 5846 8431 5910
rect 11994 5846 12041 5910
rect 12105 5846 12111 5910
rect 954 1224 1121 1288
rect 1185 1224 1191 1288
rect 4634 1224 4801 1288
rect 4865 1224 4871 1288
rect 8314 1224 8481 1288
rect 8545 1224 8551 1288
rect 11994 1224 12161 1288
rect 12225 1224 12231 1288
<< via3 >>
rect 9051 12654 9349 12752
rect 13931 12484 14229 12582
rect 6571 12314 6869 12412
rect 1691 12144 1989 12242
rect 2291 11974 2589 12072
rect 9651 11804 9949 11902
rect 341 11464 579 11732
rect 4021 11728 4259 11732
rect 4021 11468 4074 11728
rect 4074 11468 4259 11728
rect 4021 11464 4259 11468
rect 7701 11464 7939 11732
rect 11381 11464 11619 11732
rect 13331 11294 13629 11392
rect 5971 11124 6269 11222
rect 2891 10954 3189 11052
rect 5371 10784 5669 10882
rect 12731 10704 13029 10712
rect 12731 10622 12928 10704
rect 12928 10622 13029 10704
rect 12731 10614 13029 10622
rect 10251 10444 10549 10542
rect 2291 6147 2589 6545
rect 5971 6147 6269 6545
rect 9651 6147 9949 6545
rect 13331 6147 13629 6545
rect 1001 5846 1065 5910
rect 4681 5846 4745 5910
rect 8361 5846 8425 5910
rect 12041 5846 12105 5910
rect 2891 1525 3189 1923
rect 6571 1525 6869 1923
rect 10251 1525 10549 1923
rect 13931 1525 14229 1923
rect 1121 1224 1185 1288
rect 4801 1224 4865 1288
rect 8481 1224 8545 1288
rect 12161 1224 12225 1288
<< metal4 >>
rect 20 10198 260 12998
rect 340 11732 580 12998
rect 340 11464 341 11732
rect 579 11464 580 11732
rect 340 10198 580 11464
rect 660 10198 900 12998
rect 1690 12242 1990 12243
rect 1690 12144 1691 12242
rect 1989 12144 1990 12242
rect 1690 7846 1990 12144
rect 2290 12072 2590 12073
rect 2290 11974 2291 12072
rect 2589 11974 2590 12072
rect 1000 5910 1066 5911
rect 1000 5846 1001 5910
rect 1065 5846 1066 5910
rect 20 5576 260 5846
rect 340 5576 580 5846
rect 660 5576 900 5846
rect 1000 5845 1066 5846
rect 20 1136 260 1224
rect 340 1136 580 1224
rect 660 -48 900 1224
rect 1000 1140 1060 5845
rect 1690 3224 1990 7446
rect 2290 6545 2590 11974
rect 2290 6147 2291 6545
rect 2589 6147 2590 6545
rect 2290 6146 2590 6147
rect 2890 11052 3190 11053
rect 2890 10954 2891 11052
rect 3189 10954 3190 11052
rect 2890 1923 3190 10954
rect 3700 10198 3940 12998
rect 4020 11732 4260 12998
rect 4020 11464 4021 11732
rect 4259 11464 4260 11732
rect 4020 10198 4260 11464
rect 4340 10198 4580 12998
rect 6570 12412 6870 12413
rect 6570 12314 6571 12412
rect 6869 12314 6870 12412
rect 5970 11222 6270 11223
rect 5970 11124 5971 11222
rect 6269 11124 6270 11222
rect 5370 10882 5670 10883
rect 5370 10784 5371 10882
rect 5669 10784 5670 10882
rect 5370 7846 5670 10784
rect 4680 5910 4746 5911
rect 4680 5846 4681 5910
rect 4745 5846 4746 5910
rect 3700 5576 3940 5846
rect 4020 5576 4260 5846
rect 4340 5576 4580 5846
rect 4680 5845 4746 5846
rect 2890 1525 2891 1923
rect 3189 1525 3190 1923
rect 2890 1524 3190 1525
rect 1120 1288 1186 1289
rect 1120 1224 1121 1288
rect 1185 1224 1186 1288
rect 1120 1221 1186 1224
rect 1120 1140 1180 1221
rect 3700 1136 3940 1224
rect 4020 1136 4260 1224
rect 4340 -48 4580 1224
rect 4680 1140 4740 5845
rect 5370 3224 5670 7446
rect 5970 6545 6270 11124
rect 5970 6147 5971 6545
rect 6269 6147 6270 6545
rect 5970 6146 6270 6147
rect 6570 1923 6870 12314
rect 7380 10198 7620 12998
rect 7700 11732 7940 12998
rect 7700 11464 7701 11732
rect 7939 11464 7940 11732
rect 7700 10198 7940 11464
rect 8020 10198 8260 12998
rect 9050 12752 9950 12998
rect 9050 12654 9051 12752
rect 9349 12698 9950 12752
rect 9349 12654 9350 12698
rect 9050 7846 9350 12654
rect 9650 11902 9950 11903
rect 9650 11804 9651 11902
rect 9949 11804 9950 11902
rect 8360 5910 8426 5911
rect 8360 5846 8361 5910
rect 8425 5846 8426 5910
rect 7380 5576 7620 5846
rect 7700 5576 7940 5846
rect 8020 5576 8260 5846
rect 8360 5845 8426 5846
rect 6570 1525 6571 1923
rect 6869 1525 6870 1923
rect 6570 1524 6870 1525
rect 4800 1288 4866 1289
rect 4800 1224 4801 1288
rect 4865 1224 4866 1288
rect 4800 1221 4866 1224
rect 4800 1140 4860 1221
rect 7380 1136 7620 1224
rect 7700 1136 7940 1224
rect 8020 -48 8260 1224
rect 8360 1140 8420 5845
rect 9050 3224 9350 7446
rect 9650 6545 9950 11804
rect 9650 6147 9651 6545
rect 9949 6147 9950 6545
rect 9650 6146 9950 6147
rect 10250 10542 10550 10543
rect 10250 10444 10251 10542
rect 10549 10444 10550 10542
rect 10250 1923 10550 10444
rect 11060 10198 11300 12998
rect 11380 11732 11620 12998
rect 11380 11464 11381 11732
rect 11619 11464 11620 11732
rect 11380 10198 11620 11464
rect 11700 10198 11940 12998
rect 12730 12698 13630 12998
rect 12730 10712 13030 12698
rect 13930 12582 14230 12583
rect 13930 12484 13931 12582
rect 14229 12484 14230 12582
rect 12730 10614 12731 10712
rect 13029 10614 13030 10712
rect 12730 7846 13030 10614
rect 13330 11392 13630 11393
rect 13330 11294 13331 11392
rect 13629 11294 13630 11392
rect 12040 5910 12106 5911
rect 12040 5846 12041 5910
rect 12105 5846 12106 5910
rect 11060 5576 11300 5846
rect 11380 5576 11620 5846
rect 11700 5576 11940 5846
rect 12040 5845 12106 5846
rect 10250 1525 10251 1923
rect 10549 1525 10550 1923
rect 10250 1524 10550 1525
rect 8480 1288 8546 1289
rect 8480 1224 8481 1288
rect 8545 1224 8546 1288
rect 8480 1221 8546 1224
rect 8480 1140 8540 1221
rect 11060 1136 11300 1224
rect 11380 1136 11620 1224
rect 11700 -48 11940 1224
rect 12040 1140 12100 5845
rect 12730 3224 13030 7446
rect 13330 6545 13630 11294
rect 13330 6147 13331 6545
rect 13629 6147 13630 6545
rect 13330 6146 13630 6147
rect 13930 1923 14230 12484
rect 13930 1525 13931 1923
rect 14229 1525 14230 1923
rect 13930 1524 14230 1525
rect 12160 1288 12226 1289
rect 12160 1224 12161 1288
rect 12225 1224 12226 1288
rect 12160 1221 12226 1224
rect 12160 1140 12220 1221
use dev_ctrl_b2  dev_ctrl_b2_0
timestamp 1756064790
transform 1 0 11040 0 1 0
box -38 -48 3758 1140
use dev_ctrl_e2  dev_ctrl_e2_0
timestamp 1756064830
transform 1 0 0 0 1 0
box -38 -48 6868 1140
use dev_ctrl_m2  dev_ctrl_m2_0
timestamp 1756064830
transform 1 0 3680 0 1 0
box -38 -48 6868 1140
use dev_ctrl_m2  dev_ctrl_m2_1
timestamp 1756064830
transform 1 0 7360 0 1 0
box -38 -48 6868 1140
use sky130_fd_pr__nfet_g5v0d10v5_HWW8U4  sky130_fd_pr__nfet_g5v0d10v5_HWW8U4_0
timestamp 1756064685
transform 1 0 7360 0 1 11599
box -6909 -758 6909 758
use tt_asw_3v3  tt_asw_3v3_1
array 0 3 3680 0 1 -4622
timestamp 1756064685
transform 1 0 0 0 -1 5576
box 0 0 3680 4352
<< end >>
