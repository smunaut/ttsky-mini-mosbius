magic
tech sky130A
magscale 1 2
timestamp 1755863614
<< nwell >>
rect -9001 -1047 9001 1047
<< mvpmos >>
rect -8743 -750 -8543 750
rect -8485 -750 -8285 750
rect -8227 -750 -8027 750
rect -7969 -750 -7769 750
rect -7711 -750 -7511 750
rect -7453 -750 -7253 750
rect -7195 -750 -6995 750
rect -6937 -750 -6737 750
rect -6679 -750 -6479 750
rect -6421 -750 -6221 750
rect -6163 -750 -5963 750
rect -5905 -750 -5705 750
rect -5647 -750 -5447 750
rect -5389 -750 -5189 750
rect -5131 -750 -4931 750
rect -4873 -750 -4673 750
rect -4615 -750 -4415 750
rect -4357 -750 -4157 750
rect -4099 -750 -3899 750
rect -3841 -750 -3641 750
rect -3583 -750 -3383 750
rect -3325 -750 -3125 750
rect -3067 -750 -2867 750
rect -2809 -750 -2609 750
rect -2551 -750 -2351 750
rect -2293 -750 -2093 750
rect -2035 -750 -1835 750
rect -1777 -750 -1577 750
rect -1519 -750 -1319 750
rect -1261 -750 -1061 750
rect -1003 -750 -803 750
rect -745 -750 -545 750
rect -487 -750 -287 750
rect -229 -750 -29 750
rect 29 -750 229 750
rect 287 -750 487 750
rect 545 -750 745 750
rect 803 -750 1003 750
rect 1061 -750 1261 750
rect 1319 -750 1519 750
rect 1577 -750 1777 750
rect 1835 -750 2035 750
rect 2093 -750 2293 750
rect 2351 -750 2551 750
rect 2609 -750 2809 750
rect 2867 -750 3067 750
rect 3125 -750 3325 750
rect 3383 -750 3583 750
rect 3641 -750 3841 750
rect 3899 -750 4099 750
rect 4157 -750 4357 750
rect 4415 -750 4615 750
rect 4673 -750 4873 750
rect 4931 -750 5131 750
rect 5189 -750 5389 750
rect 5447 -750 5647 750
rect 5705 -750 5905 750
rect 5963 -750 6163 750
rect 6221 -750 6421 750
rect 6479 -750 6679 750
rect 6737 -750 6937 750
rect 6995 -750 7195 750
rect 7253 -750 7453 750
rect 7511 -750 7711 750
rect 7769 -750 7969 750
rect 8027 -750 8227 750
rect 8285 -750 8485 750
rect 8543 -750 8743 750
<< mvpdiff >>
rect -8801 738 -8743 750
rect -8801 -738 -8789 738
rect -8755 -738 -8743 738
rect -8801 -750 -8743 -738
rect -8543 738 -8485 750
rect -8543 -738 -8531 738
rect -8497 -738 -8485 738
rect -8543 -750 -8485 -738
rect -8285 738 -8227 750
rect -8285 -738 -8273 738
rect -8239 -738 -8227 738
rect -8285 -750 -8227 -738
rect -8027 738 -7969 750
rect -8027 -738 -8015 738
rect -7981 -738 -7969 738
rect -8027 -750 -7969 -738
rect -7769 738 -7711 750
rect -7769 -738 -7757 738
rect -7723 -738 -7711 738
rect -7769 -750 -7711 -738
rect -7511 738 -7453 750
rect -7511 -738 -7499 738
rect -7465 -738 -7453 738
rect -7511 -750 -7453 -738
rect -7253 738 -7195 750
rect -7253 -738 -7241 738
rect -7207 -738 -7195 738
rect -7253 -750 -7195 -738
rect -6995 738 -6937 750
rect -6995 -738 -6983 738
rect -6949 -738 -6937 738
rect -6995 -750 -6937 -738
rect -6737 738 -6679 750
rect -6737 -738 -6725 738
rect -6691 -738 -6679 738
rect -6737 -750 -6679 -738
rect -6479 738 -6421 750
rect -6479 -738 -6467 738
rect -6433 -738 -6421 738
rect -6479 -750 -6421 -738
rect -6221 738 -6163 750
rect -6221 -738 -6209 738
rect -6175 -738 -6163 738
rect -6221 -750 -6163 -738
rect -5963 738 -5905 750
rect -5963 -738 -5951 738
rect -5917 -738 -5905 738
rect -5963 -750 -5905 -738
rect -5705 738 -5647 750
rect -5705 -738 -5693 738
rect -5659 -738 -5647 738
rect -5705 -750 -5647 -738
rect -5447 738 -5389 750
rect -5447 -738 -5435 738
rect -5401 -738 -5389 738
rect -5447 -750 -5389 -738
rect -5189 738 -5131 750
rect -5189 -738 -5177 738
rect -5143 -738 -5131 738
rect -5189 -750 -5131 -738
rect -4931 738 -4873 750
rect -4931 -738 -4919 738
rect -4885 -738 -4873 738
rect -4931 -750 -4873 -738
rect -4673 738 -4615 750
rect -4673 -738 -4661 738
rect -4627 -738 -4615 738
rect -4673 -750 -4615 -738
rect -4415 738 -4357 750
rect -4415 -738 -4403 738
rect -4369 -738 -4357 738
rect -4415 -750 -4357 -738
rect -4157 738 -4099 750
rect -4157 -738 -4145 738
rect -4111 -738 -4099 738
rect -4157 -750 -4099 -738
rect -3899 738 -3841 750
rect -3899 -738 -3887 738
rect -3853 -738 -3841 738
rect -3899 -750 -3841 -738
rect -3641 738 -3583 750
rect -3641 -738 -3629 738
rect -3595 -738 -3583 738
rect -3641 -750 -3583 -738
rect -3383 738 -3325 750
rect -3383 -738 -3371 738
rect -3337 -738 -3325 738
rect -3383 -750 -3325 -738
rect -3125 738 -3067 750
rect -3125 -738 -3113 738
rect -3079 -738 -3067 738
rect -3125 -750 -3067 -738
rect -2867 738 -2809 750
rect -2867 -738 -2855 738
rect -2821 -738 -2809 738
rect -2867 -750 -2809 -738
rect -2609 738 -2551 750
rect -2609 -738 -2597 738
rect -2563 -738 -2551 738
rect -2609 -750 -2551 -738
rect -2351 738 -2293 750
rect -2351 -738 -2339 738
rect -2305 -738 -2293 738
rect -2351 -750 -2293 -738
rect -2093 738 -2035 750
rect -2093 -738 -2081 738
rect -2047 -738 -2035 738
rect -2093 -750 -2035 -738
rect -1835 738 -1777 750
rect -1835 -738 -1823 738
rect -1789 -738 -1777 738
rect -1835 -750 -1777 -738
rect -1577 738 -1519 750
rect -1577 -738 -1565 738
rect -1531 -738 -1519 738
rect -1577 -750 -1519 -738
rect -1319 738 -1261 750
rect -1319 -738 -1307 738
rect -1273 -738 -1261 738
rect -1319 -750 -1261 -738
rect -1061 738 -1003 750
rect -1061 -738 -1049 738
rect -1015 -738 -1003 738
rect -1061 -750 -1003 -738
rect -803 738 -745 750
rect -803 -738 -791 738
rect -757 -738 -745 738
rect -803 -750 -745 -738
rect -545 738 -487 750
rect -545 -738 -533 738
rect -499 -738 -487 738
rect -545 -750 -487 -738
rect -287 738 -229 750
rect -287 -738 -275 738
rect -241 -738 -229 738
rect -287 -750 -229 -738
rect -29 738 29 750
rect -29 -738 -17 738
rect 17 -738 29 738
rect -29 -750 29 -738
rect 229 738 287 750
rect 229 -738 241 738
rect 275 -738 287 738
rect 229 -750 287 -738
rect 487 738 545 750
rect 487 -738 499 738
rect 533 -738 545 738
rect 487 -750 545 -738
rect 745 738 803 750
rect 745 -738 757 738
rect 791 -738 803 738
rect 745 -750 803 -738
rect 1003 738 1061 750
rect 1003 -738 1015 738
rect 1049 -738 1061 738
rect 1003 -750 1061 -738
rect 1261 738 1319 750
rect 1261 -738 1273 738
rect 1307 -738 1319 738
rect 1261 -750 1319 -738
rect 1519 738 1577 750
rect 1519 -738 1531 738
rect 1565 -738 1577 738
rect 1519 -750 1577 -738
rect 1777 738 1835 750
rect 1777 -738 1789 738
rect 1823 -738 1835 738
rect 1777 -750 1835 -738
rect 2035 738 2093 750
rect 2035 -738 2047 738
rect 2081 -738 2093 738
rect 2035 -750 2093 -738
rect 2293 738 2351 750
rect 2293 -738 2305 738
rect 2339 -738 2351 738
rect 2293 -750 2351 -738
rect 2551 738 2609 750
rect 2551 -738 2563 738
rect 2597 -738 2609 738
rect 2551 -750 2609 -738
rect 2809 738 2867 750
rect 2809 -738 2821 738
rect 2855 -738 2867 738
rect 2809 -750 2867 -738
rect 3067 738 3125 750
rect 3067 -738 3079 738
rect 3113 -738 3125 738
rect 3067 -750 3125 -738
rect 3325 738 3383 750
rect 3325 -738 3337 738
rect 3371 -738 3383 738
rect 3325 -750 3383 -738
rect 3583 738 3641 750
rect 3583 -738 3595 738
rect 3629 -738 3641 738
rect 3583 -750 3641 -738
rect 3841 738 3899 750
rect 3841 -738 3853 738
rect 3887 -738 3899 738
rect 3841 -750 3899 -738
rect 4099 738 4157 750
rect 4099 -738 4111 738
rect 4145 -738 4157 738
rect 4099 -750 4157 -738
rect 4357 738 4415 750
rect 4357 -738 4369 738
rect 4403 -738 4415 738
rect 4357 -750 4415 -738
rect 4615 738 4673 750
rect 4615 -738 4627 738
rect 4661 -738 4673 738
rect 4615 -750 4673 -738
rect 4873 738 4931 750
rect 4873 -738 4885 738
rect 4919 -738 4931 738
rect 4873 -750 4931 -738
rect 5131 738 5189 750
rect 5131 -738 5143 738
rect 5177 -738 5189 738
rect 5131 -750 5189 -738
rect 5389 738 5447 750
rect 5389 -738 5401 738
rect 5435 -738 5447 738
rect 5389 -750 5447 -738
rect 5647 738 5705 750
rect 5647 -738 5659 738
rect 5693 -738 5705 738
rect 5647 -750 5705 -738
rect 5905 738 5963 750
rect 5905 -738 5917 738
rect 5951 -738 5963 738
rect 5905 -750 5963 -738
rect 6163 738 6221 750
rect 6163 -738 6175 738
rect 6209 -738 6221 738
rect 6163 -750 6221 -738
rect 6421 738 6479 750
rect 6421 -738 6433 738
rect 6467 -738 6479 738
rect 6421 -750 6479 -738
rect 6679 738 6737 750
rect 6679 -738 6691 738
rect 6725 -738 6737 738
rect 6679 -750 6737 -738
rect 6937 738 6995 750
rect 6937 -738 6949 738
rect 6983 -738 6995 738
rect 6937 -750 6995 -738
rect 7195 738 7253 750
rect 7195 -738 7207 738
rect 7241 -738 7253 738
rect 7195 -750 7253 -738
rect 7453 738 7511 750
rect 7453 -738 7465 738
rect 7499 -738 7511 738
rect 7453 -750 7511 -738
rect 7711 738 7769 750
rect 7711 -738 7723 738
rect 7757 -738 7769 738
rect 7711 -750 7769 -738
rect 7969 738 8027 750
rect 7969 -738 7981 738
rect 8015 -738 8027 738
rect 7969 -750 8027 -738
rect 8227 738 8285 750
rect 8227 -738 8239 738
rect 8273 -738 8285 738
rect 8227 -750 8285 -738
rect 8485 738 8543 750
rect 8485 -738 8497 738
rect 8531 -738 8543 738
rect 8485 -750 8543 -738
rect 8743 738 8801 750
rect 8743 -738 8755 738
rect 8789 -738 8801 738
rect 8743 -750 8801 -738
<< mvpdiffc >>
rect -8789 -738 -8755 738
rect -8531 -738 -8497 738
rect -8273 -738 -8239 738
rect -8015 -738 -7981 738
rect -7757 -738 -7723 738
rect -7499 -738 -7465 738
rect -7241 -738 -7207 738
rect -6983 -738 -6949 738
rect -6725 -738 -6691 738
rect -6467 -738 -6433 738
rect -6209 -738 -6175 738
rect -5951 -738 -5917 738
rect -5693 -738 -5659 738
rect -5435 -738 -5401 738
rect -5177 -738 -5143 738
rect -4919 -738 -4885 738
rect -4661 -738 -4627 738
rect -4403 -738 -4369 738
rect -4145 -738 -4111 738
rect -3887 -738 -3853 738
rect -3629 -738 -3595 738
rect -3371 -738 -3337 738
rect -3113 -738 -3079 738
rect -2855 -738 -2821 738
rect -2597 -738 -2563 738
rect -2339 -738 -2305 738
rect -2081 -738 -2047 738
rect -1823 -738 -1789 738
rect -1565 -738 -1531 738
rect -1307 -738 -1273 738
rect -1049 -738 -1015 738
rect -791 -738 -757 738
rect -533 -738 -499 738
rect -275 -738 -241 738
rect -17 -738 17 738
rect 241 -738 275 738
rect 499 -738 533 738
rect 757 -738 791 738
rect 1015 -738 1049 738
rect 1273 -738 1307 738
rect 1531 -738 1565 738
rect 1789 -738 1823 738
rect 2047 -738 2081 738
rect 2305 -738 2339 738
rect 2563 -738 2597 738
rect 2821 -738 2855 738
rect 3079 -738 3113 738
rect 3337 -738 3371 738
rect 3595 -738 3629 738
rect 3853 -738 3887 738
rect 4111 -738 4145 738
rect 4369 -738 4403 738
rect 4627 -738 4661 738
rect 4885 -738 4919 738
rect 5143 -738 5177 738
rect 5401 -738 5435 738
rect 5659 -738 5693 738
rect 5917 -738 5951 738
rect 6175 -738 6209 738
rect 6433 -738 6467 738
rect 6691 -738 6725 738
rect 6949 -738 6983 738
rect 7207 -738 7241 738
rect 7465 -738 7499 738
rect 7723 -738 7757 738
rect 7981 -738 8015 738
rect 8239 -738 8273 738
rect 8497 -738 8531 738
rect 8755 -738 8789 738
<< mvnsubdiff >>
rect -8935 969 8935 981
rect -8935 935 -8827 969
rect 8827 935 8935 969
rect -8935 923 8935 935
rect -8935 873 -8877 923
rect -8935 -873 -8923 873
rect -8889 -873 -8877 873
rect 8877 873 8935 923
rect -8935 -923 -8877 -873
rect 8877 -873 8889 873
rect 8923 -873 8935 873
rect 8877 -923 8935 -873
rect -8935 -935 8935 -923
rect -8935 -969 -8827 -935
rect 8827 -969 8935 -935
rect -8935 -981 8935 -969
<< mvnsubdiffcont >>
rect -8827 935 8827 969
rect -8923 -873 -8889 873
rect 8889 -873 8923 873
rect -8827 -969 8827 -935
<< poly >>
rect -8743 831 -8543 847
rect -8743 797 -8727 831
rect -8559 797 -8543 831
rect -8743 750 -8543 797
rect -8485 831 -8285 847
rect -8485 797 -8469 831
rect -8301 797 -8285 831
rect -8485 750 -8285 797
rect -8227 831 -8027 847
rect -8227 797 -8211 831
rect -8043 797 -8027 831
rect -8227 750 -8027 797
rect -7969 831 -7769 847
rect -7969 797 -7953 831
rect -7785 797 -7769 831
rect -7969 750 -7769 797
rect -7711 831 -7511 847
rect -7711 797 -7695 831
rect -7527 797 -7511 831
rect -7711 750 -7511 797
rect -7453 831 -7253 847
rect -7453 797 -7437 831
rect -7269 797 -7253 831
rect -7453 750 -7253 797
rect -7195 831 -6995 847
rect -7195 797 -7179 831
rect -7011 797 -6995 831
rect -7195 750 -6995 797
rect -6937 831 -6737 847
rect -6937 797 -6921 831
rect -6753 797 -6737 831
rect -6937 750 -6737 797
rect -6679 831 -6479 847
rect -6679 797 -6663 831
rect -6495 797 -6479 831
rect -6679 750 -6479 797
rect -6421 831 -6221 847
rect -6421 797 -6405 831
rect -6237 797 -6221 831
rect -6421 750 -6221 797
rect -6163 831 -5963 847
rect -6163 797 -6147 831
rect -5979 797 -5963 831
rect -6163 750 -5963 797
rect -5905 831 -5705 847
rect -5905 797 -5889 831
rect -5721 797 -5705 831
rect -5905 750 -5705 797
rect -5647 831 -5447 847
rect -5647 797 -5631 831
rect -5463 797 -5447 831
rect -5647 750 -5447 797
rect -5389 831 -5189 847
rect -5389 797 -5373 831
rect -5205 797 -5189 831
rect -5389 750 -5189 797
rect -5131 831 -4931 847
rect -5131 797 -5115 831
rect -4947 797 -4931 831
rect -5131 750 -4931 797
rect -4873 831 -4673 847
rect -4873 797 -4857 831
rect -4689 797 -4673 831
rect -4873 750 -4673 797
rect -4615 831 -4415 847
rect -4615 797 -4599 831
rect -4431 797 -4415 831
rect -4615 750 -4415 797
rect -4357 831 -4157 847
rect -4357 797 -4341 831
rect -4173 797 -4157 831
rect -4357 750 -4157 797
rect -4099 831 -3899 847
rect -4099 797 -4083 831
rect -3915 797 -3899 831
rect -4099 750 -3899 797
rect -3841 831 -3641 847
rect -3841 797 -3825 831
rect -3657 797 -3641 831
rect -3841 750 -3641 797
rect -3583 831 -3383 847
rect -3583 797 -3567 831
rect -3399 797 -3383 831
rect -3583 750 -3383 797
rect -3325 831 -3125 847
rect -3325 797 -3309 831
rect -3141 797 -3125 831
rect -3325 750 -3125 797
rect -3067 831 -2867 847
rect -3067 797 -3051 831
rect -2883 797 -2867 831
rect -3067 750 -2867 797
rect -2809 831 -2609 847
rect -2809 797 -2793 831
rect -2625 797 -2609 831
rect -2809 750 -2609 797
rect -2551 831 -2351 847
rect -2551 797 -2535 831
rect -2367 797 -2351 831
rect -2551 750 -2351 797
rect -2293 831 -2093 847
rect -2293 797 -2277 831
rect -2109 797 -2093 831
rect -2293 750 -2093 797
rect -2035 831 -1835 847
rect -2035 797 -2019 831
rect -1851 797 -1835 831
rect -2035 750 -1835 797
rect -1777 831 -1577 847
rect -1777 797 -1761 831
rect -1593 797 -1577 831
rect -1777 750 -1577 797
rect -1519 831 -1319 847
rect -1519 797 -1503 831
rect -1335 797 -1319 831
rect -1519 750 -1319 797
rect -1261 831 -1061 847
rect -1261 797 -1245 831
rect -1077 797 -1061 831
rect -1261 750 -1061 797
rect -1003 831 -803 847
rect -1003 797 -987 831
rect -819 797 -803 831
rect -1003 750 -803 797
rect -745 831 -545 847
rect -745 797 -729 831
rect -561 797 -545 831
rect -745 750 -545 797
rect -487 831 -287 847
rect -487 797 -471 831
rect -303 797 -287 831
rect -487 750 -287 797
rect -229 831 -29 847
rect -229 797 -213 831
rect -45 797 -29 831
rect -229 750 -29 797
rect 29 831 229 847
rect 29 797 45 831
rect 213 797 229 831
rect 29 750 229 797
rect 287 831 487 847
rect 287 797 303 831
rect 471 797 487 831
rect 287 750 487 797
rect 545 831 745 847
rect 545 797 561 831
rect 729 797 745 831
rect 545 750 745 797
rect 803 831 1003 847
rect 803 797 819 831
rect 987 797 1003 831
rect 803 750 1003 797
rect 1061 831 1261 847
rect 1061 797 1077 831
rect 1245 797 1261 831
rect 1061 750 1261 797
rect 1319 831 1519 847
rect 1319 797 1335 831
rect 1503 797 1519 831
rect 1319 750 1519 797
rect 1577 831 1777 847
rect 1577 797 1593 831
rect 1761 797 1777 831
rect 1577 750 1777 797
rect 1835 831 2035 847
rect 1835 797 1851 831
rect 2019 797 2035 831
rect 1835 750 2035 797
rect 2093 831 2293 847
rect 2093 797 2109 831
rect 2277 797 2293 831
rect 2093 750 2293 797
rect 2351 831 2551 847
rect 2351 797 2367 831
rect 2535 797 2551 831
rect 2351 750 2551 797
rect 2609 831 2809 847
rect 2609 797 2625 831
rect 2793 797 2809 831
rect 2609 750 2809 797
rect 2867 831 3067 847
rect 2867 797 2883 831
rect 3051 797 3067 831
rect 2867 750 3067 797
rect 3125 831 3325 847
rect 3125 797 3141 831
rect 3309 797 3325 831
rect 3125 750 3325 797
rect 3383 831 3583 847
rect 3383 797 3399 831
rect 3567 797 3583 831
rect 3383 750 3583 797
rect 3641 831 3841 847
rect 3641 797 3657 831
rect 3825 797 3841 831
rect 3641 750 3841 797
rect 3899 831 4099 847
rect 3899 797 3915 831
rect 4083 797 4099 831
rect 3899 750 4099 797
rect 4157 831 4357 847
rect 4157 797 4173 831
rect 4341 797 4357 831
rect 4157 750 4357 797
rect 4415 831 4615 847
rect 4415 797 4431 831
rect 4599 797 4615 831
rect 4415 750 4615 797
rect 4673 831 4873 847
rect 4673 797 4689 831
rect 4857 797 4873 831
rect 4673 750 4873 797
rect 4931 831 5131 847
rect 4931 797 4947 831
rect 5115 797 5131 831
rect 4931 750 5131 797
rect 5189 831 5389 847
rect 5189 797 5205 831
rect 5373 797 5389 831
rect 5189 750 5389 797
rect 5447 831 5647 847
rect 5447 797 5463 831
rect 5631 797 5647 831
rect 5447 750 5647 797
rect 5705 831 5905 847
rect 5705 797 5721 831
rect 5889 797 5905 831
rect 5705 750 5905 797
rect 5963 831 6163 847
rect 5963 797 5979 831
rect 6147 797 6163 831
rect 5963 750 6163 797
rect 6221 831 6421 847
rect 6221 797 6237 831
rect 6405 797 6421 831
rect 6221 750 6421 797
rect 6479 831 6679 847
rect 6479 797 6495 831
rect 6663 797 6679 831
rect 6479 750 6679 797
rect 6737 831 6937 847
rect 6737 797 6753 831
rect 6921 797 6937 831
rect 6737 750 6937 797
rect 6995 831 7195 847
rect 6995 797 7011 831
rect 7179 797 7195 831
rect 6995 750 7195 797
rect 7253 831 7453 847
rect 7253 797 7269 831
rect 7437 797 7453 831
rect 7253 750 7453 797
rect 7511 831 7711 847
rect 7511 797 7527 831
rect 7695 797 7711 831
rect 7511 750 7711 797
rect 7769 831 7969 847
rect 7769 797 7785 831
rect 7953 797 7969 831
rect 7769 750 7969 797
rect 8027 831 8227 847
rect 8027 797 8043 831
rect 8211 797 8227 831
rect 8027 750 8227 797
rect 8285 831 8485 847
rect 8285 797 8301 831
rect 8469 797 8485 831
rect 8285 750 8485 797
rect 8543 831 8743 847
rect 8543 797 8559 831
rect 8727 797 8743 831
rect 8543 750 8743 797
rect -8743 -797 -8543 -750
rect -8743 -831 -8727 -797
rect -8559 -831 -8543 -797
rect -8743 -847 -8543 -831
rect -8485 -797 -8285 -750
rect -8485 -831 -8469 -797
rect -8301 -831 -8285 -797
rect -8485 -847 -8285 -831
rect -8227 -797 -8027 -750
rect -8227 -831 -8211 -797
rect -8043 -831 -8027 -797
rect -8227 -847 -8027 -831
rect -7969 -797 -7769 -750
rect -7969 -831 -7953 -797
rect -7785 -831 -7769 -797
rect -7969 -847 -7769 -831
rect -7711 -797 -7511 -750
rect -7711 -831 -7695 -797
rect -7527 -831 -7511 -797
rect -7711 -847 -7511 -831
rect -7453 -797 -7253 -750
rect -7453 -831 -7437 -797
rect -7269 -831 -7253 -797
rect -7453 -847 -7253 -831
rect -7195 -797 -6995 -750
rect -7195 -831 -7179 -797
rect -7011 -831 -6995 -797
rect -7195 -847 -6995 -831
rect -6937 -797 -6737 -750
rect -6937 -831 -6921 -797
rect -6753 -831 -6737 -797
rect -6937 -847 -6737 -831
rect -6679 -797 -6479 -750
rect -6679 -831 -6663 -797
rect -6495 -831 -6479 -797
rect -6679 -847 -6479 -831
rect -6421 -797 -6221 -750
rect -6421 -831 -6405 -797
rect -6237 -831 -6221 -797
rect -6421 -847 -6221 -831
rect -6163 -797 -5963 -750
rect -6163 -831 -6147 -797
rect -5979 -831 -5963 -797
rect -6163 -847 -5963 -831
rect -5905 -797 -5705 -750
rect -5905 -831 -5889 -797
rect -5721 -831 -5705 -797
rect -5905 -847 -5705 -831
rect -5647 -797 -5447 -750
rect -5647 -831 -5631 -797
rect -5463 -831 -5447 -797
rect -5647 -847 -5447 -831
rect -5389 -797 -5189 -750
rect -5389 -831 -5373 -797
rect -5205 -831 -5189 -797
rect -5389 -847 -5189 -831
rect -5131 -797 -4931 -750
rect -5131 -831 -5115 -797
rect -4947 -831 -4931 -797
rect -5131 -847 -4931 -831
rect -4873 -797 -4673 -750
rect -4873 -831 -4857 -797
rect -4689 -831 -4673 -797
rect -4873 -847 -4673 -831
rect -4615 -797 -4415 -750
rect -4615 -831 -4599 -797
rect -4431 -831 -4415 -797
rect -4615 -847 -4415 -831
rect -4357 -797 -4157 -750
rect -4357 -831 -4341 -797
rect -4173 -831 -4157 -797
rect -4357 -847 -4157 -831
rect -4099 -797 -3899 -750
rect -4099 -831 -4083 -797
rect -3915 -831 -3899 -797
rect -4099 -847 -3899 -831
rect -3841 -797 -3641 -750
rect -3841 -831 -3825 -797
rect -3657 -831 -3641 -797
rect -3841 -847 -3641 -831
rect -3583 -797 -3383 -750
rect -3583 -831 -3567 -797
rect -3399 -831 -3383 -797
rect -3583 -847 -3383 -831
rect -3325 -797 -3125 -750
rect -3325 -831 -3309 -797
rect -3141 -831 -3125 -797
rect -3325 -847 -3125 -831
rect -3067 -797 -2867 -750
rect -3067 -831 -3051 -797
rect -2883 -831 -2867 -797
rect -3067 -847 -2867 -831
rect -2809 -797 -2609 -750
rect -2809 -831 -2793 -797
rect -2625 -831 -2609 -797
rect -2809 -847 -2609 -831
rect -2551 -797 -2351 -750
rect -2551 -831 -2535 -797
rect -2367 -831 -2351 -797
rect -2551 -847 -2351 -831
rect -2293 -797 -2093 -750
rect -2293 -831 -2277 -797
rect -2109 -831 -2093 -797
rect -2293 -847 -2093 -831
rect -2035 -797 -1835 -750
rect -2035 -831 -2019 -797
rect -1851 -831 -1835 -797
rect -2035 -847 -1835 -831
rect -1777 -797 -1577 -750
rect -1777 -831 -1761 -797
rect -1593 -831 -1577 -797
rect -1777 -847 -1577 -831
rect -1519 -797 -1319 -750
rect -1519 -831 -1503 -797
rect -1335 -831 -1319 -797
rect -1519 -847 -1319 -831
rect -1261 -797 -1061 -750
rect -1261 -831 -1245 -797
rect -1077 -831 -1061 -797
rect -1261 -847 -1061 -831
rect -1003 -797 -803 -750
rect -1003 -831 -987 -797
rect -819 -831 -803 -797
rect -1003 -847 -803 -831
rect -745 -797 -545 -750
rect -745 -831 -729 -797
rect -561 -831 -545 -797
rect -745 -847 -545 -831
rect -487 -797 -287 -750
rect -487 -831 -471 -797
rect -303 -831 -287 -797
rect -487 -847 -287 -831
rect -229 -797 -29 -750
rect -229 -831 -213 -797
rect -45 -831 -29 -797
rect -229 -847 -29 -831
rect 29 -797 229 -750
rect 29 -831 45 -797
rect 213 -831 229 -797
rect 29 -847 229 -831
rect 287 -797 487 -750
rect 287 -831 303 -797
rect 471 -831 487 -797
rect 287 -847 487 -831
rect 545 -797 745 -750
rect 545 -831 561 -797
rect 729 -831 745 -797
rect 545 -847 745 -831
rect 803 -797 1003 -750
rect 803 -831 819 -797
rect 987 -831 1003 -797
rect 803 -847 1003 -831
rect 1061 -797 1261 -750
rect 1061 -831 1077 -797
rect 1245 -831 1261 -797
rect 1061 -847 1261 -831
rect 1319 -797 1519 -750
rect 1319 -831 1335 -797
rect 1503 -831 1519 -797
rect 1319 -847 1519 -831
rect 1577 -797 1777 -750
rect 1577 -831 1593 -797
rect 1761 -831 1777 -797
rect 1577 -847 1777 -831
rect 1835 -797 2035 -750
rect 1835 -831 1851 -797
rect 2019 -831 2035 -797
rect 1835 -847 2035 -831
rect 2093 -797 2293 -750
rect 2093 -831 2109 -797
rect 2277 -831 2293 -797
rect 2093 -847 2293 -831
rect 2351 -797 2551 -750
rect 2351 -831 2367 -797
rect 2535 -831 2551 -797
rect 2351 -847 2551 -831
rect 2609 -797 2809 -750
rect 2609 -831 2625 -797
rect 2793 -831 2809 -797
rect 2609 -847 2809 -831
rect 2867 -797 3067 -750
rect 2867 -831 2883 -797
rect 3051 -831 3067 -797
rect 2867 -847 3067 -831
rect 3125 -797 3325 -750
rect 3125 -831 3141 -797
rect 3309 -831 3325 -797
rect 3125 -847 3325 -831
rect 3383 -797 3583 -750
rect 3383 -831 3399 -797
rect 3567 -831 3583 -797
rect 3383 -847 3583 -831
rect 3641 -797 3841 -750
rect 3641 -831 3657 -797
rect 3825 -831 3841 -797
rect 3641 -847 3841 -831
rect 3899 -797 4099 -750
rect 3899 -831 3915 -797
rect 4083 -831 4099 -797
rect 3899 -847 4099 -831
rect 4157 -797 4357 -750
rect 4157 -831 4173 -797
rect 4341 -831 4357 -797
rect 4157 -847 4357 -831
rect 4415 -797 4615 -750
rect 4415 -831 4431 -797
rect 4599 -831 4615 -797
rect 4415 -847 4615 -831
rect 4673 -797 4873 -750
rect 4673 -831 4689 -797
rect 4857 -831 4873 -797
rect 4673 -847 4873 -831
rect 4931 -797 5131 -750
rect 4931 -831 4947 -797
rect 5115 -831 5131 -797
rect 4931 -847 5131 -831
rect 5189 -797 5389 -750
rect 5189 -831 5205 -797
rect 5373 -831 5389 -797
rect 5189 -847 5389 -831
rect 5447 -797 5647 -750
rect 5447 -831 5463 -797
rect 5631 -831 5647 -797
rect 5447 -847 5647 -831
rect 5705 -797 5905 -750
rect 5705 -831 5721 -797
rect 5889 -831 5905 -797
rect 5705 -847 5905 -831
rect 5963 -797 6163 -750
rect 5963 -831 5979 -797
rect 6147 -831 6163 -797
rect 5963 -847 6163 -831
rect 6221 -797 6421 -750
rect 6221 -831 6237 -797
rect 6405 -831 6421 -797
rect 6221 -847 6421 -831
rect 6479 -797 6679 -750
rect 6479 -831 6495 -797
rect 6663 -831 6679 -797
rect 6479 -847 6679 -831
rect 6737 -797 6937 -750
rect 6737 -831 6753 -797
rect 6921 -831 6937 -797
rect 6737 -847 6937 -831
rect 6995 -797 7195 -750
rect 6995 -831 7011 -797
rect 7179 -831 7195 -797
rect 6995 -847 7195 -831
rect 7253 -797 7453 -750
rect 7253 -831 7269 -797
rect 7437 -831 7453 -797
rect 7253 -847 7453 -831
rect 7511 -797 7711 -750
rect 7511 -831 7527 -797
rect 7695 -831 7711 -797
rect 7511 -847 7711 -831
rect 7769 -797 7969 -750
rect 7769 -831 7785 -797
rect 7953 -831 7969 -797
rect 7769 -847 7969 -831
rect 8027 -797 8227 -750
rect 8027 -831 8043 -797
rect 8211 -831 8227 -797
rect 8027 -847 8227 -831
rect 8285 -797 8485 -750
rect 8285 -831 8301 -797
rect 8469 -831 8485 -797
rect 8285 -847 8485 -831
rect 8543 -797 8743 -750
rect 8543 -831 8559 -797
rect 8727 -831 8743 -797
rect 8543 -847 8743 -831
<< polycont >>
rect -8727 797 -8559 831
rect -8469 797 -8301 831
rect -8211 797 -8043 831
rect -7953 797 -7785 831
rect -7695 797 -7527 831
rect -7437 797 -7269 831
rect -7179 797 -7011 831
rect -6921 797 -6753 831
rect -6663 797 -6495 831
rect -6405 797 -6237 831
rect -6147 797 -5979 831
rect -5889 797 -5721 831
rect -5631 797 -5463 831
rect -5373 797 -5205 831
rect -5115 797 -4947 831
rect -4857 797 -4689 831
rect -4599 797 -4431 831
rect -4341 797 -4173 831
rect -4083 797 -3915 831
rect -3825 797 -3657 831
rect -3567 797 -3399 831
rect -3309 797 -3141 831
rect -3051 797 -2883 831
rect -2793 797 -2625 831
rect -2535 797 -2367 831
rect -2277 797 -2109 831
rect -2019 797 -1851 831
rect -1761 797 -1593 831
rect -1503 797 -1335 831
rect -1245 797 -1077 831
rect -987 797 -819 831
rect -729 797 -561 831
rect -471 797 -303 831
rect -213 797 -45 831
rect 45 797 213 831
rect 303 797 471 831
rect 561 797 729 831
rect 819 797 987 831
rect 1077 797 1245 831
rect 1335 797 1503 831
rect 1593 797 1761 831
rect 1851 797 2019 831
rect 2109 797 2277 831
rect 2367 797 2535 831
rect 2625 797 2793 831
rect 2883 797 3051 831
rect 3141 797 3309 831
rect 3399 797 3567 831
rect 3657 797 3825 831
rect 3915 797 4083 831
rect 4173 797 4341 831
rect 4431 797 4599 831
rect 4689 797 4857 831
rect 4947 797 5115 831
rect 5205 797 5373 831
rect 5463 797 5631 831
rect 5721 797 5889 831
rect 5979 797 6147 831
rect 6237 797 6405 831
rect 6495 797 6663 831
rect 6753 797 6921 831
rect 7011 797 7179 831
rect 7269 797 7437 831
rect 7527 797 7695 831
rect 7785 797 7953 831
rect 8043 797 8211 831
rect 8301 797 8469 831
rect 8559 797 8727 831
rect -8727 -831 -8559 -797
rect -8469 -831 -8301 -797
rect -8211 -831 -8043 -797
rect -7953 -831 -7785 -797
rect -7695 -831 -7527 -797
rect -7437 -831 -7269 -797
rect -7179 -831 -7011 -797
rect -6921 -831 -6753 -797
rect -6663 -831 -6495 -797
rect -6405 -831 -6237 -797
rect -6147 -831 -5979 -797
rect -5889 -831 -5721 -797
rect -5631 -831 -5463 -797
rect -5373 -831 -5205 -797
rect -5115 -831 -4947 -797
rect -4857 -831 -4689 -797
rect -4599 -831 -4431 -797
rect -4341 -831 -4173 -797
rect -4083 -831 -3915 -797
rect -3825 -831 -3657 -797
rect -3567 -831 -3399 -797
rect -3309 -831 -3141 -797
rect -3051 -831 -2883 -797
rect -2793 -831 -2625 -797
rect -2535 -831 -2367 -797
rect -2277 -831 -2109 -797
rect -2019 -831 -1851 -797
rect -1761 -831 -1593 -797
rect -1503 -831 -1335 -797
rect -1245 -831 -1077 -797
rect -987 -831 -819 -797
rect -729 -831 -561 -797
rect -471 -831 -303 -797
rect -213 -831 -45 -797
rect 45 -831 213 -797
rect 303 -831 471 -797
rect 561 -831 729 -797
rect 819 -831 987 -797
rect 1077 -831 1245 -797
rect 1335 -831 1503 -797
rect 1593 -831 1761 -797
rect 1851 -831 2019 -797
rect 2109 -831 2277 -797
rect 2367 -831 2535 -797
rect 2625 -831 2793 -797
rect 2883 -831 3051 -797
rect 3141 -831 3309 -797
rect 3399 -831 3567 -797
rect 3657 -831 3825 -797
rect 3915 -831 4083 -797
rect 4173 -831 4341 -797
rect 4431 -831 4599 -797
rect 4689 -831 4857 -797
rect 4947 -831 5115 -797
rect 5205 -831 5373 -797
rect 5463 -831 5631 -797
rect 5721 -831 5889 -797
rect 5979 -831 6147 -797
rect 6237 -831 6405 -797
rect 6495 -831 6663 -797
rect 6753 -831 6921 -797
rect 7011 -831 7179 -797
rect 7269 -831 7437 -797
rect 7527 -831 7695 -797
rect 7785 -831 7953 -797
rect 8043 -831 8211 -797
rect 8301 -831 8469 -797
rect 8559 -831 8727 -797
<< locali >>
rect -8923 935 -8827 969
rect 8827 935 8923 969
rect -8923 873 -8889 935
rect 8889 873 8923 935
rect -8743 797 -8727 831
rect -8559 797 -8543 831
rect -8485 797 -8469 831
rect -8301 797 -8285 831
rect -8227 797 -8211 831
rect -8043 797 -8027 831
rect -7969 797 -7953 831
rect -7785 797 -7769 831
rect -7711 797 -7695 831
rect -7527 797 -7511 831
rect -7453 797 -7437 831
rect -7269 797 -7253 831
rect -7195 797 -7179 831
rect -7011 797 -6995 831
rect -6937 797 -6921 831
rect -6753 797 -6737 831
rect -6679 797 -6663 831
rect -6495 797 -6479 831
rect -6421 797 -6405 831
rect -6237 797 -6221 831
rect -6163 797 -6147 831
rect -5979 797 -5963 831
rect -5905 797 -5889 831
rect -5721 797 -5705 831
rect -5647 797 -5631 831
rect -5463 797 -5447 831
rect -5389 797 -5373 831
rect -5205 797 -5189 831
rect -5131 797 -5115 831
rect -4947 797 -4931 831
rect -4873 797 -4857 831
rect -4689 797 -4673 831
rect -4615 797 -4599 831
rect -4431 797 -4415 831
rect -4357 797 -4341 831
rect -4173 797 -4157 831
rect -4099 797 -4083 831
rect -3915 797 -3899 831
rect -3841 797 -3825 831
rect -3657 797 -3641 831
rect -3583 797 -3567 831
rect -3399 797 -3383 831
rect -3325 797 -3309 831
rect -3141 797 -3125 831
rect -3067 797 -3051 831
rect -2883 797 -2867 831
rect -2809 797 -2793 831
rect -2625 797 -2609 831
rect -2551 797 -2535 831
rect -2367 797 -2351 831
rect -2293 797 -2277 831
rect -2109 797 -2093 831
rect -2035 797 -2019 831
rect -1851 797 -1835 831
rect -1777 797 -1761 831
rect -1593 797 -1577 831
rect -1519 797 -1503 831
rect -1335 797 -1319 831
rect -1261 797 -1245 831
rect -1077 797 -1061 831
rect -1003 797 -987 831
rect -819 797 -803 831
rect -745 797 -729 831
rect -561 797 -545 831
rect -487 797 -471 831
rect -303 797 -287 831
rect -229 797 -213 831
rect -45 797 -29 831
rect 29 797 45 831
rect 213 797 229 831
rect 287 797 303 831
rect 471 797 487 831
rect 545 797 561 831
rect 729 797 745 831
rect 803 797 819 831
rect 987 797 1003 831
rect 1061 797 1077 831
rect 1245 797 1261 831
rect 1319 797 1335 831
rect 1503 797 1519 831
rect 1577 797 1593 831
rect 1761 797 1777 831
rect 1835 797 1851 831
rect 2019 797 2035 831
rect 2093 797 2109 831
rect 2277 797 2293 831
rect 2351 797 2367 831
rect 2535 797 2551 831
rect 2609 797 2625 831
rect 2793 797 2809 831
rect 2867 797 2883 831
rect 3051 797 3067 831
rect 3125 797 3141 831
rect 3309 797 3325 831
rect 3383 797 3399 831
rect 3567 797 3583 831
rect 3641 797 3657 831
rect 3825 797 3841 831
rect 3899 797 3915 831
rect 4083 797 4099 831
rect 4157 797 4173 831
rect 4341 797 4357 831
rect 4415 797 4431 831
rect 4599 797 4615 831
rect 4673 797 4689 831
rect 4857 797 4873 831
rect 4931 797 4947 831
rect 5115 797 5131 831
rect 5189 797 5205 831
rect 5373 797 5389 831
rect 5447 797 5463 831
rect 5631 797 5647 831
rect 5705 797 5721 831
rect 5889 797 5905 831
rect 5963 797 5979 831
rect 6147 797 6163 831
rect 6221 797 6237 831
rect 6405 797 6421 831
rect 6479 797 6495 831
rect 6663 797 6679 831
rect 6737 797 6753 831
rect 6921 797 6937 831
rect 6995 797 7011 831
rect 7179 797 7195 831
rect 7253 797 7269 831
rect 7437 797 7453 831
rect 7511 797 7527 831
rect 7695 797 7711 831
rect 7769 797 7785 831
rect 7953 797 7969 831
rect 8027 797 8043 831
rect 8211 797 8227 831
rect 8285 797 8301 831
rect 8469 797 8485 831
rect 8543 797 8559 831
rect 8727 797 8743 831
rect -8789 738 -8755 754
rect -8789 -754 -8755 -738
rect -8531 738 -8497 754
rect -8531 -754 -8497 -738
rect -8273 738 -8239 754
rect -8273 -754 -8239 -738
rect -8015 738 -7981 754
rect -8015 -754 -7981 -738
rect -7757 738 -7723 754
rect -7757 -754 -7723 -738
rect -7499 738 -7465 754
rect -7499 -754 -7465 -738
rect -7241 738 -7207 754
rect -7241 -754 -7207 -738
rect -6983 738 -6949 754
rect -6983 -754 -6949 -738
rect -6725 738 -6691 754
rect -6725 -754 -6691 -738
rect -6467 738 -6433 754
rect -6467 -754 -6433 -738
rect -6209 738 -6175 754
rect -6209 -754 -6175 -738
rect -5951 738 -5917 754
rect -5951 -754 -5917 -738
rect -5693 738 -5659 754
rect -5693 -754 -5659 -738
rect -5435 738 -5401 754
rect -5435 -754 -5401 -738
rect -5177 738 -5143 754
rect -5177 -754 -5143 -738
rect -4919 738 -4885 754
rect -4919 -754 -4885 -738
rect -4661 738 -4627 754
rect -4661 -754 -4627 -738
rect -4403 738 -4369 754
rect -4403 -754 -4369 -738
rect -4145 738 -4111 754
rect -4145 -754 -4111 -738
rect -3887 738 -3853 754
rect -3887 -754 -3853 -738
rect -3629 738 -3595 754
rect -3629 -754 -3595 -738
rect -3371 738 -3337 754
rect -3371 -754 -3337 -738
rect -3113 738 -3079 754
rect -3113 -754 -3079 -738
rect -2855 738 -2821 754
rect -2855 -754 -2821 -738
rect -2597 738 -2563 754
rect -2597 -754 -2563 -738
rect -2339 738 -2305 754
rect -2339 -754 -2305 -738
rect -2081 738 -2047 754
rect -2081 -754 -2047 -738
rect -1823 738 -1789 754
rect -1823 -754 -1789 -738
rect -1565 738 -1531 754
rect -1565 -754 -1531 -738
rect -1307 738 -1273 754
rect -1307 -754 -1273 -738
rect -1049 738 -1015 754
rect -1049 -754 -1015 -738
rect -791 738 -757 754
rect -791 -754 -757 -738
rect -533 738 -499 754
rect -533 -754 -499 -738
rect -275 738 -241 754
rect -275 -754 -241 -738
rect -17 738 17 754
rect -17 -754 17 -738
rect 241 738 275 754
rect 241 -754 275 -738
rect 499 738 533 754
rect 499 -754 533 -738
rect 757 738 791 754
rect 757 -754 791 -738
rect 1015 738 1049 754
rect 1015 -754 1049 -738
rect 1273 738 1307 754
rect 1273 -754 1307 -738
rect 1531 738 1565 754
rect 1531 -754 1565 -738
rect 1789 738 1823 754
rect 1789 -754 1823 -738
rect 2047 738 2081 754
rect 2047 -754 2081 -738
rect 2305 738 2339 754
rect 2305 -754 2339 -738
rect 2563 738 2597 754
rect 2563 -754 2597 -738
rect 2821 738 2855 754
rect 2821 -754 2855 -738
rect 3079 738 3113 754
rect 3079 -754 3113 -738
rect 3337 738 3371 754
rect 3337 -754 3371 -738
rect 3595 738 3629 754
rect 3595 -754 3629 -738
rect 3853 738 3887 754
rect 3853 -754 3887 -738
rect 4111 738 4145 754
rect 4111 -754 4145 -738
rect 4369 738 4403 754
rect 4369 -754 4403 -738
rect 4627 738 4661 754
rect 4627 -754 4661 -738
rect 4885 738 4919 754
rect 4885 -754 4919 -738
rect 5143 738 5177 754
rect 5143 -754 5177 -738
rect 5401 738 5435 754
rect 5401 -754 5435 -738
rect 5659 738 5693 754
rect 5659 -754 5693 -738
rect 5917 738 5951 754
rect 5917 -754 5951 -738
rect 6175 738 6209 754
rect 6175 -754 6209 -738
rect 6433 738 6467 754
rect 6433 -754 6467 -738
rect 6691 738 6725 754
rect 6691 -754 6725 -738
rect 6949 738 6983 754
rect 6949 -754 6983 -738
rect 7207 738 7241 754
rect 7207 -754 7241 -738
rect 7465 738 7499 754
rect 7465 -754 7499 -738
rect 7723 738 7757 754
rect 7723 -754 7757 -738
rect 7981 738 8015 754
rect 7981 -754 8015 -738
rect 8239 738 8273 754
rect 8239 -754 8273 -738
rect 8497 738 8531 754
rect 8497 -754 8531 -738
rect 8755 738 8789 754
rect 8755 -754 8789 -738
rect -8743 -831 -8727 -797
rect -8559 -831 -8543 -797
rect -8485 -831 -8469 -797
rect -8301 -831 -8285 -797
rect -8227 -831 -8211 -797
rect -8043 -831 -8027 -797
rect -7969 -831 -7953 -797
rect -7785 -831 -7769 -797
rect -7711 -831 -7695 -797
rect -7527 -831 -7511 -797
rect -7453 -831 -7437 -797
rect -7269 -831 -7253 -797
rect -7195 -831 -7179 -797
rect -7011 -831 -6995 -797
rect -6937 -831 -6921 -797
rect -6753 -831 -6737 -797
rect -6679 -831 -6663 -797
rect -6495 -831 -6479 -797
rect -6421 -831 -6405 -797
rect -6237 -831 -6221 -797
rect -6163 -831 -6147 -797
rect -5979 -831 -5963 -797
rect -5905 -831 -5889 -797
rect -5721 -831 -5705 -797
rect -5647 -831 -5631 -797
rect -5463 -831 -5447 -797
rect -5389 -831 -5373 -797
rect -5205 -831 -5189 -797
rect -5131 -831 -5115 -797
rect -4947 -831 -4931 -797
rect -4873 -831 -4857 -797
rect -4689 -831 -4673 -797
rect -4615 -831 -4599 -797
rect -4431 -831 -4415 -797
rect -4357 -831 -4341 -797
rect -4173 -831 -4157 -797
rect -4099 -831 -4083 -797
rect -3915 -831 -3899 -797
rect -3841 -831 -3825 -797
rect -3657 -831 -3641 -797
rect -3583 -831 -3567 -797
rect -3399 -831 -3383 -797
rect -3325 -831 -3309 -797
rect -3141 -831 -3125 -797
rect -3067 -831 -3051 -797
rect -2883 -831 -2867 -797
rect -2809 -831 -2793 -797
rect -2625 -831 -2609 -797
rect -2551 -831 -2535 -797
rect -2367 -831 -2351 -797
rect -2293 -831 -2277 -797
rect -2109 -831 -2093 -797
rect -2035 -831 -2019 -797
rect -1851 -831 -1835 -797
rect -1777 -831 -1761 -797
rect -1593 -831 -1577 -797
rect -1519 -831 -1503 -797
rect -1335 -831 -1319 -797
rect -1261 -831 -1245 -797
rect -1077 -831 -1061 -797
rect -1003 -831 -987 -797
rect -819 -831 -803 -797
rect -745 -831 -729 -797
rect -561 -831 -545 -797
rect -487 -831 -471 -797
rect -303 -831 -287 -797
rect -229 -831 -213 -797
rect -45 -831 -29 -797
rect 29 -831 45 -797
rect 213 -831 229 -797
rect 287 -831 303 -797
rect 471 -831 487 -797
rect 545 -831 561 -797
rect 729 -831 745 -797
rect 803 -831 819 -797
rect 987 -831 1003 -797
rect 1061 -831 1077 -797
rect 1245 -831 1261 -797
rect 1319 -831 1335 -797
rect 1503 -831 1519 -797
rect 1577 -831 1593 -797
rect 1761 -831 1777 -797
rect 1835 -831 1851 -797
rect 2019 -831 2035 -797
rect 2093 -831 2109 -797
rect 2277 -831 2293 -797
rect 2351 -831 2367 -797
rect 2535 -831 2551 -797
rect 2609 -831 2625 -797
rect 2793 -831 2809 -797
rect 2867 -831 2883 -797
rect 3051 -831 3067 -797
rect 3125 -831 3141 -797
rect 3309 -831 3325 -797
rect 3383 -831 3399 -797
rect 3567 -831 3583 -797
rect 3641 -831 3657 -797
rect 3825 -831 3841 -797
rect 3899 -831 3915 -797
rect 4083 -831 4099 -797
rect 4157 -831 4173 -797
rect 4341 -831 4357 -797
rect 4415 -831 4431 -797
rect 4599 -831 4615 -797
rect 4673 -831 4689 -797
rect 4857 -831 4873 -797
rect 4931 -831 4947 -797
rect 5115 -831 5131 -797
rect 5189 -831 5205 -797
rect 5373 -831 5389 -797
rect 5447 -831 5463 -797
rect 5631 -831 5647 -797
rect 5705 -831 5721 -797
rect 5889 -831 5905 -797
rect 5963 -831 5979 -797
rect 6147 -831 6163 -797
rect 6221 -831 6237 -797
rect 6405 -831 6421 -797
rect 6479 -831 6495 -797
rect 6663 -831 6679 -797
rect 6737 -831 6753 -797
rect 6921 -831 6937 -797
rect 6995 -831 7011 -797
rect 7179 -831 7195 -797
rect 7253 -831 7269 -797
rect 7437 -831 7453 -797
rect 7511 -831 7527 -797
rect 7695 -831 7711 -797
rect 7769 -831 7785 -797
rect 7953 -831 7969 -797
rect 8027 -831 8043 -797
rect 8211 -831 8227 -797
rect 8285 -831 8301 -797
rect 8469 -831 8485 -797
rect 8543 -831 8559 -797
rect 8727 -831 8743 -797
rect -8923 -935 -8889 -873
rect 8889 -935 8923 -873
rect -8923 -969 -8827 -935
rect 8827 -969 8923 -935
<< viali >>
rect -8727 797 -8559 831
rect -8469 797 -8301 831
rect -8211 797 -8043 831
rect -7953 797 -7785 831
rect -7695 797 -7527 831
rect -7437 797 -7269 831
rect -7179 797 -7011 831
rect -6921 797 -6753 831
rect -6663 797 -6495 831
rect -6405 797 -6237 831
rect -6147 797 -5979 831
rect -5889 797 -5721 831
rect -5631 797 -5463 831
rect -5373 797 -5205 831
rect -5115 797 -4947 831
rect -4857 797 -4689 831
rect -4599 797 -4431 831
rect -4341 797 -4173 831
rect -4083 797 -3915 831
rect -3825 797 -3657 831
rect -3567 797 -3399 831
rect -3309 797 -3141 831
rect -3051 797 -2883 831
rect -2793 797 -2625 831
rect -2535 797 -2367 831
rect -2277 797 -2109 831
rect -2019 797 -1851 831
rect -1761 797 -1593 831
rect -1503 797 -1335 831
rect -1245 797 -1077 831
rect -987 797 -819 831
rect -729 797 -561 831
rect -471 797 -303 831
rect -213 797 -45 831
rect 45 797 213 831
rect 303 797 471 831
rect 561 797 729 831
rect 819 797 987 831
rect 1077 797 1245 831
rect 1335 797 1503 831
rect 1593 797 1761 831
rect 1851 797 2019 831
rect 2109 797 2277 831
rect 2367 797 2535 831
rect 2625 797 2793 831
rect 2883 797 3051 831
rect 3141 797 3309 831
rect 3399 797 3567 831
rect 3657 797 3825 831
rect 3915 797 4083 831
rect 4173 797 4341 831
rect 4431 797 4599 831
rect 4689 797 4857 831
rect 4947 797 5115 831
rect 5205 797 5373 831
rect 5463 797 5631 831
rect 5721 797 5889 831
rect 5979 797 6147 831
rect 6237 797 6405 831
rect 6495 797 6663 831
rect 6753 797 6921 831
rect 7011 797 7179 831
rect 7269 797 7437 831
rect 7527 797 7695 831
rect 7785 797 7953 831
rect 8043 797 8211 831
rect 8301 797 8469 831
rect 8559 797 8727 831
rect -8789 -738 -8755 738
rect -8531 -738 -8497 738
rect -8273 -738 -8239 738
rect -8015 -738 -7981 738
rect -7757 -738 -7723 738
rect -7499 -738 -7465 738
rect -7241 -738 -7207 738
rect -6983 -738 -6949 738
rect -6725 -738 -6691 738
rect -6467 -738 -6433 738
rect -6209 -738 -6175 738
rect -5951 -738 -5917 738
rect -5693 -738 -5659 738
rect -5435 -738 -5401 738
rect -5177 -738 -5143 738
rect -4919 -738 -4885 738
rect -4661 -738 -4627 738
rect -4403 -738 -4369 738
rect -4145 -738 -4111 738
rect -3887 -738 -3853 738
rect -3629 -738 -3595 738
rect -3371 -738 -3337 738
rect -3113 -738 -3079 738
rect -2855 -738 -2821 738
rect -2597 -738 -2563 738
rect -2339 -738 -2305 738
rect -2081 -738 -2047 738
rect -1823 -738 -1789 738
rect -1565 -738 -1531 738
rect -1307 -738 -1273 738
rect -1049 -738 -1015 738
rect -791 -738 -757 738
rect -533 -738 -499 738
rect -275 -738 -241 738
rect -17 -738 17 738
rect 241 -738 275 738
rect 499 -738 533 738
rect 757 -738 791 738
rect 1015 -738 1049 738
rect 1273 -738 1307 738
rect 1531 -738 1565 738
rect 1789 -738 1823 738
rect 2047 -738 2081 738
rect 2305 -738 2339 738
rect 2563 -738 2597 738
rect 2821 -738 2855 738
rect 3079 -738 3113 738
rect 3337 -738 3371 738
rect 3595 -738 3629 738
rect 3853 -738 3887 738
rect 4111 -738 4145 738
rect 4369 -738 4403 738
rect 4627 -738 4661 738
rect 4885 -738 4919 738
rect 5143 -738 5177 738
rect 5401 -738 5435 738
rect 5659 -738 5693 738
rect 5917 -738 5951 738
rect 6175 -738 6209 738
rect 6433 -738 6467 738
rect 6691 -738 6725 738
rect 6949 -738 6983 738
rect 7207 -738 7241 738
rect 7465 -738 7499 738
rect 7723 -738 7757 738
rect 7981 -738 8015 738
rect 8239 -738 8273 738
rect 8497 -738 8531 738
rect 8755 -738 8789 738
rect -8727 -831 -8559 -797
rect -8469 -831 -8301 -797
rect -8211 -831 -8043 -797
rect -7953 -831 -7785 -797
rect -7695 -831 -7527 -797
rect -7437 -831 -7269 -797
rect -7179 -831 -7011 -797
rect -6921 -831 -6753 -797
rect -6663 -831 -6495 -797
rect -6405 -831 -6237 -797
rect -6147 -831 -5979 -797
rect -5889 -831 -5721 -797
rect -5631 -831 -5463 -797
rect -5373 -831 -5205 -797
rect -5115 -831 -4947 -797
rect -4857 -831 -4689 -797
rect -4599 -831 -4431 -797
rect -4341 -831 -4173 -797
rect -4083 -831 -3915 -797
rect -3825 -831 -3657 -797
rect -3567 -831 -3399 -797
rect -3309 -831 -3141 -797
rect -3051 -831 -2883 -797
rect -2793 -831 -2625 -797
rect -2535 -831 -2367 -797
rect -2277 -831 -2109 -797
rect -2019 -831 -1851 -797
rect -1761 -831 -1593 -797
rect -1503 -831 -1335 -797
rect -1245 -831 -1077 -797
rect -987 -831 -819 -797
rect -729 -831 -561 -797
rect -471 -831 -303 -797
rect -213 -831 -45 -797
rect 45 -831 213 -797
rect 303 -831 471 -797
rect 561 -831 729 -797
rect 819 -831 987 -797
rect 1077 -831 1245 -797
rect 1335 -831 1503 -797
rect 1593 -831 1761 -797
rect 1851 -831 2019 -797
rect 2109 -831 2277 -797
rect 2367 -831 2535 -797
rect 2625 -831 2793 -797
rect 2883 -831 3051 -797
rect 3141 -831 3309 -797
rect 3399 -831 3567 -797
rect 3657 -831 3825 -797
rect 3915 -831 4083 -797
rect 4173 -831 4341 -797
rect 4431 -831 4599 -797
rect 4689 -831 4857 -797
rect 4947 -831 5115 -797
rect 5205 -831 5373 -797
rect 5463 -831 5631 -797
rect 5721 -831 5889 -797
rect 5979 -831 6147 -797
rect 6237 -831 6405 -797
rect 6495 -831 6663 -797
rect 6753 -831 6921 -797
rect 7011 -831 7179 -797
rect 7269 -831 7437 -797
rect 7527 -831 7695 -797
rect 7785 -831 7953 -797
rect 8043 -831 8211 -797
rect 8301 -831 8469 -797
rect 8559 -831 8727 -797
<< metal1 >>
rect -8739 831 -8547 837
rect -8739 797 -8727 831
rect -8559 797 -8547 831
rect -8739 791 -8547 797
rect -8481 831 -8289 837
rect -8481 797 -8469 831
rect -8301 797 -8289 831
rect -8481 791 -8289 797
rect -8223 831 -8031 837
rect -8223 797 -8211 831
rect -8043 797 -8031 831
rect -8223 791 -8031 797
rect -7965 831 -7773 837
rect -7965 797 -7953 831
rect -7785 797 -7773 831
rect -7965 791 -7773 797
rect -7707 831 -7515 837
rect -7707 797 -7695 831
rect -7527 797 -7515 831
rect -7707 791 -7515 797
rect -7449 831 -7257 837
rect -7449 797 -7437 831
rect -7269 797 -7257 831
rect -7449 791 -7257 797
rect -7191 831 -6999 837
rect -7191 797 -7179 831
rect -7011 797 -6999 831
rect -7191 791 -6999 797
rect -6933 831 -6741 837
rect -6933 797 -6921 831
rect -6753 797 -6741 831
rect -6933 791 -6741 797
rect -6675 831 -6483 837
rect -6675 797 -6663 831
rect -6495 797 -6483 831
rect -6675 791 -6483 797
rect -6417 831 -6225 837
rect -6417 797 -6405 831
rect -6237 797 -6225 831
rect -6417 791 -6225 797
rect -6159 831 -5967 837
rect -6159 797 -6147 831
rect -5979 797 -5967 831
rect -6159 791 -5967 797
rect -5901 831 -5709 837
rect -5901 797 -5889 831
rect -5721 797 -5709 831
rect -5901 791 -5709 797
rect -5643 831 -5451 837
rect -5643 797 -5631 831
rect -5463 797 -5451 831
rect -5643 791 -5451 797
rect -5385 831 -5193 837
rect -5385 797 -5373 831
rect -5205 797 -5193 831
rect -5385 791 -5193 797
rect -5127 831 -4935 837
rect -5127 797 -5115 831
rect -4947 797 -4935 831
rect -5127 791 -4935 797
rect -4869 831 -4677 837
rect -4869 797 -4857 831
rect -4689 797 -4677 831
rect -4869 791 -4677 797
rect -4611 831 -4419 837
rect -4611 797 -4599 831
rect -4431 797 -4419 831
rect -4611 791 -4419 797
rect -4353 831 -4161 837
rect -4353 797 -4341 831
rect -4173 797 -4161 831
rect -4353 791 -4161 797
rect -4095 831 -3903 837
rect -4095 797 -4083 831
rect -3915 797 -3903 831
rect -4095 791 -3903 797
rect -3837 831 -3645 837
rect -3837 797 -3825 831
rect -3657 797 -3645 831
rect -3837 791 -3645 797
rect -3579 831 -3387 837
rect -3579 797 -3567 831
rect -3399 797 -3387 831
rect -3579 791 -3387 797
rect -3321 831 -3129 837
rect -3321 797 -3309 831
rect -3141 797 -3129 831
rect -3321 791 -3129 797
rect -3063 831 -2871 837
rect -3063 797 -3051 831
rect -2883 797 -2871 831
rect -3063 791 -2871 797
rect -2805 831 -2613 837
rect -2805 797 -2793 831
rect -2625 797 -2613 831
rect -2805 791 -2613 797
rect -2547 831 -2355 837
rect -2547 797 -2535 831
rect -2367 797 -2355 831
rect -2547 791 -2355 797
rect -2289 831 -2097 837
rect -2289 797 -2277 831
rect -2109 797 -2097 831
rect -2289 791 -2097 797
rect -2031 831 -1839 837
rect -2031 797 -2019 831
rect -1851 797 -1839 831
rect -2031 791 -1839 797
rect -1773 831 -1581 837
rect -1773 797 -1761 831
rect -1593 797 -1581 831
rect -1773 791 -1581 797
rect -1515 831 -1323 837
rect -1515 797 -1503 831
rect -1335 797 -1323 831
rect -1515 791 -1323 797
rect -1257 831 -1065 837
rect -1257 797 -1245 831
rect -1077 797 -1065 831
rect -1257 791 -1065 797
rect -999 831 -807 837
rect -999 797 -987 831
rect -819 797 -807 831
rect -999 791 -807 797
rect -741 831 -549 837
rect -741 797 -729 831
rect -561 797 -549 831
rect -741 791 -549 797
rect -483 831 -291 837
rect -483 797 -471 831
rect -303 797 -291 831
rect -483 791 -291 797
rect -225 831 -33 837
rect -225 797 -213 831
rect -45 797 -33 831
rect -225 791 -33 797
rect 33 831 225 837
rect 33 797 45 831
rect 213 797 225 831
rect 33 791 225 797
rect 291 831 483 837
rect 291 797 303 831
rect 471 797 483 831
rect 291 791 483 797
rect 549 831 741 837
rect 549 797 561 831
rect 729 797 741 831
rect 549 791 741 797
rect 807 831 999 837
rect 807 797 819 831
rect 987 797 999 831
rect 807 791 999 797
rect 1065 831 1257 837
rect 1065 797 1077 831
rect 1245 797 1257 831
rect 1065 791 1257 797
rect 1323 831 1515 837
rect 1323 797 1335 831
rect 1503 797 1515 831
rect 1323 791 1515 797
rect 1581 831 1773 837
rect 1581 797 1593 831
rect 1761 797 1773 831
rect 1581 791 1773 797
rect 1839 831 2031 837
rect 1839 797 1851 831
rect 2019 797 2031 831
rect 1839 791 2031 797
rect 2097 831 2289 837
rect 2097 797 2109 831
rect 2277 797 2289 831
rect 2097 791 2289 797
rect 2355 831 2547 837
rect 2355 797 2367 831
rect 2535 797 2547 831
rect 2355 791 2547 797
rect 2613 831 2805 837
rect 2613 797 2625 831
rect 2793 797 2805 831
rect 2613 791 2805 797
rect 2871 831 3063 837
rect 2871 797 2883 831
rect 3051 797 3063 831
rect 2871 791 3063 797
rect 3129 831 3321 837
rect 3129 797 3141 831
rect 3309 797 3321 831
rect 3129 791 3321 797
rect 3387 831 3579 837
rect 3387 797 3399 831
rect 3567 797 3579 831
rect 3387 791 3579 797
rect 3645 831 3837 837
rect 3645 797 3657 831
rect 3825 797 3837 831
rect 3645 791 3837 797
rect 3903 831 4095 837
rect 3903 797 3915 831
rect 4083 797 4095 831
rect 3903 791 4095 797
rect 4161 831 4353 837
rect 4161 797 4173 831
rect 4341 797 4353 831
rect 4161 791 4353 797
rect 4419 831 4611 837
rect 4419 797 4431 831
rect 4599 797 4611 831
rect 4419 791 4611 797
rect 4677 831 4869 837
rect 4677 797 4689 831
rect 4857 797 4869 831
rect 4677 791 4869 797
rect 4935 831 5127 837
rect 4935 797 4947 831
rect 5115 797 5127 831
rect 4935 791 5127 797
rect 5193 831 5385 837
rect 5193 797 5205 831
rect 5373 797 5385 831
rect 5193 791 5385 797
rect 5451 831 5643 837
rect 5451 797 5463 831
rect 5631 797 5643 831
rect 5451 791 5643 797
rect 5709 831 5901 837
rect 5709 797 5721 831
rect 5889 797 5901 831
rect 5709 791 5901 797
rect 5967 831 6159 837
rect 5967 797 5979 831
rect 6147 797 6159 831
rect 5967 791 6159 797
rect 6225 831 6417 837
rect 6225 797 6237 831
rect 6405 797 6417 831
rect 6225 791 6417 797
rect 6483 831 6675 837
rect 6483 797 6495 831
rect 6663 797 6675 831
rect 6483 791 6675 797
rect 6741 831 6933 837
rect 6741 797 6753 831
rect 6921 797 6933 831
rect 6741 791 6933 797
rect 6999 831 7191 837
rect 6999 797 7011 831
rect 7179 797 7191 831
rect 6999 791 7191 797
rect 7257 831 7449 837
rect 7257 797 7269 831
rect 7437 797 7449 831
rect 7257 791 7449 797
rect 7515 831 7707 837
rect 7515 797 7527 831
rect 7695 797 7707 831
rect 7515 791 7707 797
rect 7773 831 7965 837
rect 7773 797 7785 831
rect 7953 797 7965 831
rect 7773 791 7965 797
rect 8031 831 8223 837
rect 8031 797 8043 831
rect 8211 797 8223 831
rect 8031 791 8223 797
rect 8289 831 8481 837
rect 8289 797 8301 831
rect 8469 797 8481 831
rect 8289 791 8481 797
rect 8547 831 8739 837
rect 8547 797 8559 831
rect 8727 797 8739 831
rect 8547 791 8739 797
rect -8795 738 -8749 750
rect -8795 -738 -8789 738
rect -8755 -738 -8749 738
rect -8795 -750 -8749 -738
rect -8537 738 -8491 750
rect -8537 -738 -8531 738
rect -8497 -738 -8491 738
rect -8537 -750 -8491 -738
rect -8279 738 -8233 750
rect -8279 -738 -8273 738
rect -8239 -738 -8233 738
rect -8279 -750 -8233 -738
rect -8021 738 -7975 750
rect -8021 -738 -8015 738
rect -7981 -738 -7975 738
rect -8021 -750 -7975 -738
rect -7763 738 -7717 750
rect -7763 -738 -7757 738
rect -7723 -738 -7717 738
rect -7763 -750 -7717 -738
rect -7505 738 -7459 750
rect -7505 -738 -7499 738
rect -7465 -738 -7459 738
rect -7505 -750 -7459 -738
rect -7247 738 -7201 750
rect -7247 -738 -7241 738
rect -7207 -738 -7201 738
rect -7247 -750 -7201 -738
rect -6989 738 -6943 750
rect -6989 -738 -6983 738
rect -6949 -738 -6943 738
rect -6989 -750 -6943 -738
rect -6731 738 -6685 750
rect -6731 -738 -6725 738
rect -6691 -738 -6685 738
rect -6731 -750 -6685 -738
rect -6473 738 -6427 750
rect -6473 -738 -6467 738
rect -6433 -738 -6427 738
rect -6473 -750 -6427 -738
rect -6215 738 -6169 750
rect -6215 -738 -6209 738
rect -6175 -738 -6169 738
rect -6215 -750 -6169 -738
rect -5957 738 -5911 750
rect -5957 -738 -5951 738
rect -5917 -738 -5911 738
rect -5957 -750 -5911 -738
rect -5699 738 -5653 750
rect -5699 -738 -5693 738
rect -5659 -738 -5653 738
rect -5699 -750 -5653 -738
rect -5441 738 -5395 750
rect -5441 -738 -5435 738
rect -5401 -738 -5395 738
rect -5441 -750 -5395 -738
rect -5183 738 -5137 750
rect -5183 -738 -5177 738
rect -5143 -738 -5137 738
rect -5183 -750 -5137 -738
rect -4925 738 -4879 750
rect -4925 -738 -4919 738
rect -4885 -738 -4879 738
rect -4925 -750 -4879 -738
rect -4667 738 -4621 750
rect -4667 -738 -4661 738
rect -4627 -738 -4621 738
rect -4667 -750 -4621 -738
rect -4409 738 -4363 750
rect -4409 -738 -4403 738
rect -4369 -738 -4363 738
rect -4409 -750 -4363 -738
rect -4151 738 -4105 750
rect -4151 -738 -4145 738
rect -4111 -738 -4105 738
rect -4151 -750 -4105 -738
rect -3893 738 -3847 750
rect -3893 -738 -3887 738
rect -3853 -738 -3847 738
rect -3893 -750 -3847 -738
rect -3635 738 -3589 750
rect -3635 -738 -3629 738
rect -3595 -738 -3589 738
rect -3635 -750 -3589 -738
rect -3377 738 -3331 750
rect -3377 -738 -3371 738
rect -3337 -738 -3331 738
rect -3377 -750 -3331 -738
rect -3119 738 -3073 750
rect -3119 -738 -3113 738
rect -3079 -738 -3073 738
rect -3119 -750 -3073 -738
rect -2861 738 -2815 750
rect -2861 -738 -2855 738
rect -2821 -738 -2815 738
rect -2861 -750 -2815 -738
rect -2603 738 -2557 750
rect -2603 -738 -2597 738
rect -2563 -738 -2557 738
rect -2603 -750 -2557 -738
rect -2345 738 -2299 750
rect -2345 -738 -2339 738
rect -2305 -738 -2299 738
rect -2345 -750 -2299 -738
rect -2087 738 -2041 750
rect -2087 -738 -2081 738
rect -2047 -738 -2041 738
rect -2087 -750 -2041 -738
rect -1829 738 -1783 750
rect -1829 -738 -1823 738
rect -1789 -738 -1783 738
rect -1829 -750 -1783 -738
rect -1571 738 -1525 750
rect -1571 -738 -1565 738
rect -1531 -738 -1525 738
rect -1571 -750 -1525 -738
rect -1313 738 -1267 750
rect -1313 -738 -1307 738
rect -1273 -738 -1267 738
rect -1313 -750 -1267 -738
rect -1055 738 -1009 750
rect -1055 -738 -1049 738
rect -1015 -738 -1009 738
rect -1055 -750 -1009 -738
rect -797 738 -751 750
rect -797 -738 -791 738
rect -757 -738 -751 738
rect -797 -750 -751 -738
rect -539 738 -493 750
rect -539 -738 -533 738
rect -499 -738 -493 738
rect -539 -750 -493 -738
rect -281 738 -235 750
rect -281 -738 -275 738
rect -241 -738 -235 738
rect -281 -750 -235 -738
rect -23 738 23 750
rect -23 -738 -17 738
rect 17 -738 23 738
rect -23 -750 23 -738
rect 235 738 281 750
rect 235 -738 241 738
rect 275 -738 281 738
rect 235 -750 281 -738
rect 493 738 539 750
rect 493 -738 499 738
rect 533 -738 539 738
rect 493 -750 539 -738
rect 751 738 797 750
rect 751 -738 757 738
rect 791 -738 797 738
rect 751 -750 797 -738
rect 1009 738 1055 750
rect 1009 -738 1015 738
rect 1049 -738 1055 738
rect 1009 -750 1055 -738
rect 1267 738 1313 750
rect 1267 -738 1273 738
rect 1307 -738 1313 738
rect 1267 -750 1313 -738
rect 1525 738 1571 750
rect 1525 -738 1531 738
rect 1565 -738 1571 738
rect 1525 -750 1571 -738
rect 1783 738 1829 750
rect 1783 -738 1789 738
rect 1823 -738 1829 738
rect 1783 -750 1829 -738
rect 2041 738 2087 750
rect 2041 -738 2047 738
rect 2081 -738 2087 738
rect 2041 -750 2087 -738
rect 2299 738 2345 750
rect 2299 -738 2305 738
rect 2339 -738 2345 738
rect 2299 -750 2345 -738
rect 2557 738 2603 750
rect 2557 -738 2563 738
rect 2597 -738 2603 738
rect 2557 -750 2603 -738
rect 2815 738 2861 750
rect 2815 -738 2821 738
rect 2855 -738 2861 738
rect 2815 -750 2861 -738
rect 3073 738 3119 750
rect 3073 -738 3079 738
rect 3113 -738 3119 738
rect 3073 -750 3119 -738
rect 3331 738 3377 750
rect 3331 -738 3337 738
rect 3371 -738 3377 738
rect 3331 -750 3377 -738
rect 3589 738 3635 750
rect 3589 -738 3595 738
rect 3629 -738 3635 738
rect 3589 -750 3635 -738
rect 3847 738 3893 750
rect 3847 -738 3853 738
rect 3887 -738 3893 738
rect 3847 -750 3893 -738
rect 4105 738 4151 750
rect 4105 -738 4111 738
rect 4145 -738 4151 738
rect 4105 -750 4151 -738
rect 4363 738 4409 750
rect 4363 -738 4369 738
rect 4403 -738 4409 738
rect 4363 -750 4409 -738
rect 4621 738 4667 750
rect 4621 -738 4627 738
rect 4661 -738 4667 738
rect 4621 -750 4667 -738
rect 4879 738 4925 750
rect 4879 -738 4885 738
rect 4919 -738 4925 738
rect 4879 -750 4925 -738
rect 5137 738 5183 750
rect 5137 -738 5143 738
rect 5177 -738 5183 738
rect 5137 -750 5183 -738
rect 5395 738 5441 750
rect 5395 -738 5401 738
rect 5435 -738 5441 738
rect 5395 -750 5441 -738
rect 5653 738 5699 750
rect 5653 -738 5659 738
rect 5693 -738 5699 738
rect 5653 -750 5699 -738
rect 5911 738 5957 750
rect 5911 -738 5917 738
rect 5951 -738 5957 738
rect 5911 -750 5957 -738
rect 6169 738 6215 750
rect 6169 -738 6175 738
rect 6209 -738 6215 738
rect 6169 -750 6215 -738
rect 6427 738 6473 750
rect 6427 -738 6433 738
rect 6467 -738 6473 738
rect 6427 -750 6473 -738
rect 6685 738 6731 750
rect 6685 -738 6691 738
rect 6725 -738 6731 738
rect 6685 -750 6731 -738
rect 6943 738 6989 750
rect 6943 -738 6949 738
rect 6983 -738 6989 738
rect 6943 -750 6989 -738
rect 7201 738 7247 750
rect 7201 -738 7207 738
rect 7241 -738 7247 738
rect 7201 -750 7247 -738
rect 7459 738 7505 750
rect 7459 -738 7465 738
rect 7499 -738 7505 738
rect 7459 -750 7505 -738
rect 7717 738 7763 750
rect 7717 -738 7723 738
rect 7757 -738 7763 738
rect 7717 -750 7763 -738
rect 7975 738 8021 750
rect 7975 -738 7981 738
rect 8015 -738 8021 738
rect 7975 -750 8021 -738
rect 8233 738 8279 750
rect 8233 -738 8239 738
rect 8273 -738 8279 738
rect 8233 -750 8279 -738
rect 8491 738 8537 750
rect 8491 -738 8497 738
rect 8531 -738 8537 738
rect 8491 -750 8537 -738
rect 8749 738 8795 750
rect 8749 -738 8755 738
rect 8789 -738 8795 738
rect 8749 -750 8795 -738
rect -8739 -797 -8547 -791
rect -8739 -831 -8727 -797
rect -8559 -831 -8547 -797
rect -8739 -837 -8547 -831
rect -8481 -797 -8289 -791
rect -8481 -831 -8469 -797
rect -8301 -831 -8289 -797
rect -8481 -837 -8289 -831
rect -8223 -797 -8031 -791
rect -8223 -831 -8211 -797
rect -8043 -831 -8031 -797
rect -8223 -837 -8031 -831
rect -7965 -797 -7773 -791
rect -7965 -831 -7953 -797
rect -7785 -831 -7773 -797
rect -7965 -837 -7773 -831
rect -7707 -797 -7515 -791
rect -7707 -831 -7695 -797
rect -7527 -831 -7515 -797
rect -7707 -837 -7515 -831
rect -7449 -797 -7257 -791
rect -7449 -831 -7437 -797
rect -7269 -831 -7257 -797
rect -7449 -837 -7257 -831
rect -7191 -797 -6999 -791
rect -7191 -831 -7179 -797
rect -7011 -831 -6999 -797
rect -7191 -837 -6999 -831
rect -6933 -797 -6741 -791
rect -6933 -831 -6921 -797
rect -6753 -831 -6741 -797
rect -6933 -837 -6741 -831
rect -6675 -797 -6483 -791
rect -6675 -831 -6663 -797
rect -6495 -831 -6483 -797
rect -6675 -837 -6483 -831
rect -6417 -797 -6225 -791
rect -6417 -831 -6405 -797
rect -6237 -831 -6225 -797
rect -6417 -837 -6225 -831
rect -6159 -797 -5967 -791
rect -6159 -831 -6147 -797
rect -5979 -831 -5967 -797
rect -6159 -837 -5967 -831
rect -5901 -797 -5709 -791
rect -5901 -831 -5889 -797
rect -5721 -831 -5709 -797
rect -5901 -837 -5709 -831
rect -5643 -797 -5451 -791
rect -5643 -831 -5631 -797
rect -5463 -831 -5451 -797
rect -5643 -837 -5451 -831
rect -5385 -797 -5193 -791
rect -5385 -831 -5373 -797
rect -5205 -831 -5193 -797
rect -5385 -837 -5193 -831
rect -5127 -797 -4935 -791
rect -5127 -831 -5115 -797
rect -4947 -831 -4935 -797
rect -5127 -837 -4935 -831
rect -4869 -797 -4677 -791
rect -4869 -831 -4857 -797
rect -4689 -831 -4677 -797
rect -4869 -837 -4677 -831
rect -4611 -797 -4419 -791
rect -4611 -831 -4599 -797
rect -4431 -831 -4419 -797
rect -4611 -837 -4419 -831
rect -4353 -797 -4161 -791
rect -4353 -831 -4341 -797
rect -4173 -831 -4161 -797
rect -4353 -837 -4161 -831
rect -4095 -797 -3903 -791
rect -4095 -831 -4083 -797
rect -3915 -831 -3903 -797
rect -4095 -837 -3903 -831
rect -3837 -797 -3645 -791
rect -3837 -831 -3825 -797
rect -3657 -831 -3645 -797
rect -3837 -837 -3645 -831
rect -3579 -797 -3387 -791
rect -3579 -831 -3567 -797
rect -3399 -831 -3387 -797
rect -3579 -837 -3387 -831
rect -3321 -797 -3129 -791
rect -3321 -831 -3309 -797
rect -3141 -831 -3129 -797
rect -3321 -837 -3129 -831
rect -3063 -797 -2871 -791
rect -3063 -831 -3051 -797
rect -2883 -831 -2871 -797
rect -3063 -837 -2871 -831
rect -2805 -797 -2613 -791
rect -2805 -831 -2793 -797
rect -2625 -831 -2613 -797
rect -2805 -837 -2613 -831
rect -2547 -797 -2355 -791
rect -2547 -831 -2535 -797
rect -2367 -831 -2355 -797
rect -2547 -837 -2355 -831
rect -2289 -797 -2097 -791
rect -2289 -831 -2277 -797
rect -2109 -831 -2097 -797
rect -2289 -837 -2097 -831
rect -2031 -797 -1839 -791
rect -2031 -831 -2019 -797
rect -1851 -831 -1839 -797
rect -2031 -837 -1839 -831
rect -1773 -797 -1581 -791
rect -1773 -831 -1761 -797
rect -1593 -831 -1581 -797
rect -1773 -837 -1581 -831
rect -1515 -797 -1323 -791
rect -1515 -831 -1503 -797
rect -1335 -831 -1323 -797
rect -1515 -837 -1323 -831
rect -1257 -797 -1065 -791
rect -1257 -831 -1245 -797
rect -1077 -831 -1065 -797
rect -1257 -837 -1065 -831
rect -999 -797 -807 -791
rect -999 -831 -987 -797
rect -819 -831 -807 -797
rect -999 -837 -807 -831
rect -741 -797 -549 -791
rect -741 -831 -729 -797
rect -561 -831 -549 -797
rect -741 -837 -549 -831
rect -483 -797 -291 -791
rect -483 -831 -471 -797
rect -303 -831 -291 -797
rect -483 -837 -291 -831
rect -225 -797 -33 -791
rect -225 -831 -213 -797
rect -45 -831 -33 -797
rect -225 -837 -33 -831
rect 33 -797 225 -791
rect 33 -831 45 -797
rect 213 -831 225 -797
rect 33 -837 225 -831
rect 291 -797 483 -791
rect 291 -831 303 -797
rect 471 -831 483 -797
rect 291 -837 483 -831
rect 549 -797 741 -791
rect 549 -831 561 -797
rect 729 -831 741 -797
rect 549 -837 741 -831
rect 807 -797 999 -791
rect 807 -831 819 -797
rect 987 -831 999 -797
rect 807 -837 999 -831
rect 1065 -797 1257 -791
rect 1065 -831 1077 -797
rect 1245 -831 1257 -797
rect 1065 -837 1257 -831
rect 1323 -797 1515 -791
rect 1323 -831 1335 -797
rect 1503 -831 1515 -797
rect 1323 -837 1515 -831
rect 1581 -797 1773 -791
rect 1581 -831 1593 -797
rect 1761 -831 1773 -797
rect 1581 -837 1773 -831
rect 1839 -797 2031 -791
rect 1839 -831 1851 -797
rect 2019 -831 2031 -797
rect 1839 -837 2031 -831
rect 2097 -797 2289 -791
rect 2097 -831 2109 -797
rect 2277 -831 2289 -797
rect 2097 -837 2289 -831
rect 2355 -797 2547 -791
rect 2355 -831 2367 -797
rect 2535 -831 2547 -797
rect 2355 -837 2547 -831
rect 2613 -797 2805 -791
rect 2613 -831 2625 -797
rect 2793 -831 2805 -797
rect 2613 -837 2805 -831
rect 2871 -797 3063 -791
rect 2871 -831 2883 -797
rect 3051 -831 3063 -797
rect 2871 -837 3063 -831
rect 3129 -797 3321 -791
rect 3129 -831 3141 -797
rect 3309 -831 3321 -797
rect 3129 -837 3321 -831
rect 3387 -797 3579 -791
rect 3387 -831 3399 -797
rect 3567 -831 3579 -797
rect 3387 -837 3579 -831
rect 3645 -797 3837 -791
rect 3645 -831 3657 -797
rect 3825 -831 3837 -797
rect 3645 -837 3837 -831
rect 3903 -797 4095 -791
rect 3903 -831 3915 -797
rect 4083 -831 4095 -797
rect 3903 -837 4095 -831
rect 4161 -797 4353 -791
rect 4161 -831 4173 -797
rect 4341 -831 4353 -797
rect 4161 -837 4353 -831
rect 4419 -797 4611 -791
rect 4419 -831 4431 -797
rect 4599 -831 4611 -797
rect 4419 -837 4611 -831
rect 4677 -797 4869 -791
rect 4677 -831 4689 -797
rect 4857 -831 4869 -797
rect 4677 -837 4869 -831
rect 4935 -797 5127 -791
rect 4935 -831 4947 -797
rect 5115 -831 5127 -797
rect 4935 -837 5127 -831
rect 5193 -797 5385 -791
rect 5193 -831 5205 -797
rect 5373 -831 5385 -797
rect 5193 -837 5385 -831
rect 5451 -797 5643 -791
rect 5451 -831 5463 -797
rect 5631 -831 5643 -797
rect 5451 -837 5643 -831
rect 5709 -797 5901 -791
rect 5709 -831 5721 -797
rect 5889 -831 5901 -797
rect 5709 -837 5901 -831
rect 5967 -797 6159 -791
rect 5967 -831 5979 -797
rect 6147 -831 6159 -797
rect 5967 -837 6159 -831
rect 6225 -797 6417 -791
rect 6225 -831 6237 -797
rect 6405 -831 6417 -797
rect 6225 -837 6417 -831
rect 6483 -797 6675 -791
rect 6483 -831 6495 -797
rect 6663 -831 6675 -797
rect 6483 -837 6675 -831
rect 6741 -797 6933 -791
rect 6741 -831 6753 -797
rect 6921 -831 6933 -797
rect 6741 -837 6933 -831
rect 6999 -797 7191 -791
rect 6999 -831 7011 -797
rect 7179 -831 7191 -797
rect 6999 -837 7191 -831
rect 7257 -797 7449 -791
rect 7257 -831 7269 -797
rect 7437 -831 7449 -797
rect 7257 -837 7449 -831
rect 7515 -797 7707 -791
rect 7515 -831 7527 -797
rect 7695 -831 7707 -797
rect 7515 -837 7707 -831
rect 7773 -797 7965 -791
rect 7773 -831 7785 -797
rect 7953 -831 7965 -797
rect 7773 -837 7965 -831
rect 8031 -797 8223 -791
rect 8031 -831 8043 -797
rect 8211 -831 8223 -797
rect 8031 -837 8223 -831
rect 8289 -797 8481 -791
rect 8289 -831 8301 -797
rect 8469 -831 8481 -797
rect 8289 -837 8481 -831
rect 8547 -797 8739 -791
rect 8547 -831 8559 -797
rect 8727 -831 8739 -797
rect 8547 -837 8739 -831
<< labels >>
rlabel mvnsubdiffcont 0 -952 0 -952 0 B
port 1 nsew
rlabel mvpdiffc -8772 0 -8772 0 0 D0
port 2 nsew
rlabel polycont -8643 814 -8643 814 0 G0
port 3 nsew
rlabel mvpdiffc -8514 0 -8514 0 0 S1
port 4 nsew
rlabel polycont -8385 814 -8385 814 0 G1
port 5 nsew
rlabel mvpdiffc -8256 0 -8256 0 0 D2
port 6 nsew
rlabel polycont -8127 814 -8127 814 0 G2
port 7 nsew
rlabel mvpdiffc -7998 0 -7998 0 0 S3
port 8 nsew
rlabel polycont -7869 814 -7869 814 0 G3
port 9 nsew
rlabel mvpdiffc -7740 0 -7740 0 0 D4
port 10 nsew
rlabel polycont -7611 814 -7611 814 0 G4
port 11 nsew
rlabel mvpdiffc -7482 0 -7482 0 0 S5
port 12 nsew
rlabel polycont -7353 814 -7353 814 0 G5
port 13 nsew
rlabel mvpdiffc -7224 0 -7224 0 0 D6
port 14 nsew
rlabel polycont -7095 814 -7095 814 0 G6
port 15 nsew
rlabel mvpdiffc -6966 0 -6966 0 0 S7
port 16 nsew
rlabel polycont -6837 814 -6837 814 0 G7
port 17 nsew
rlabel mvpdiffc -6708 0 -6708 0 0 D8
port 18 nsew
rlabel polycont -6579 814 -6579 814 0 G8
port 19 nsew
rlabel mvpdiffc -6450 0 -6450 0 0 S9
port 20 nsew
rlabel polycont -6321 814 -6321 814 0 G9
port 21 nsew
rlabel mvpdiffc -6192 0 -6192 0 0 D10
port 22 nsew
rlabel polycont -6063 814 -6063 814 0 G10
port 23 nsew
rlabel mvpdiffc -5934 0 -5934 0 0 S11
port 24 nsew
rlabel polycont -5805 814 -5805 814 0 G11
port 25 nsew
rlabel mvpdiffc -5676 0 -5676 0 0 D12
port 26 nsew
rlabel polycont -5547 814 -5547 814 0 G12
port 27 nsew
rlabel mvpdiffc -5418 0 -5418 0 0 S13
port 28 nsew
rlabel polycont -5289 814 -5289 814 0 G13
port 29 nsew
rlabel mvpdiffc -5160 0 -5160 0 0 D14
port 30 nsew
rlabel polycont -5031 814 -5031 814 0 G14
port 31 nsew
rlabel mvpdiffc -4902 0 -4902 0 0 S15
port 32 nsew
rlabel polycont -4773 814 -4773 814 0 G15
port 33 nsew
rlabel mvpdiffc -4644 0 -4644 0 0 D16
port 34 nsew
rlabel polycont -4515 814 -4515 814 0 G16
port 35 nsew
rlabel mvpdiffc -4386 0 -4386 0 0 S17
port 36 nsew
rlabel polycont -4257 814 -4257 814 0 G17
port 37 nsew
rlabel mvpdiffc -4128 0 -4128 0 0 D18
port 38 nsew
rlabel polycont -3999 814 -3999 814 0 G18
port 39 nsew
rlabel mvpdiffc -3870 0 -3870 0 0 S19
port 40 nsew
rlabel polycont -3741 814 -3741 814 0 G19
port 41 nsew
rlabel mvpdiffc -3612 0 -3612 0 0 D20
port 42 nsew
rlabel polycont -3483 814 -3483 814 0 G20
port 43 nsew
rlabel mvpdiffc -3354 0 -3354 0 0 S21
port 44 nsew
rlabel polycont -3225 814 -3225 814 0 G21
port 45 nsew
rlabel mvpdiffc -3096 0 -3096 0 0 D22
port 46 nsew
rlabel polycont -2967 814 -2967 814 0 G22
port 47 nsew
rlabel mvpdiffc -2838 0 -2838 0 0 S23
port 48 nsew
rlabel polycont -2709 814 -2709 814 0 G23
port 49 nsew
rlabel mvpdiffc -2580 0 -2580 0 0 D24
port 50 nsew
rlabel polycont -2451 814 -2451 814 0 G24
port 51 nsew
rlabel mvpdiffc -2322 0 -2322 0 0 S25
port 52 nsew
rlabel polycont -2193 814 -2193 814 0 G25
port 53 nsew
rlabel mvpdiffc -2064 0 -2064 0 0 D26
port 54 nsew
rlabel polycont -1935 814 -1935 814 0 G26
port 55 nsew
rlabel mvpdiffc -1806 0 -1806 0 0 S27
port 56 nsew
rlabel polycont -1677 814 -1677 814 0 G27
port 57 nsew
rlabel mvpdiffc -1548 0 -1548 0 0 D28
port 58 nsew
rlabel polycont -1419 814 -1419 814 0 G28
port 59 nsew
rlabel mvpdiffc -1290 0 -1290 0 0 S29
port 60 nsew
rlabel polycont -1161 814 -1161 814 0 G29
port 61 nsew
rlabel mvpdiffc -1032 0 -1032 0 0 D30
port 62 nsew
rlabel polycont -903 814 -903 814 0 G30
port 63 nsew
rlabel mvpdiffc -774 0 -774 0 0 S31
port 64 nsew
rlabel polycont -645 814 -645 814 0 G31
port 65 nsew
rlabel mvpdiffc -516 0 -516 0 0 D32
port 66 nsew
rlabel polycont -387 814 -387 814 0 G32
port 67 nsew
rlabel mvpdiffc -258 0 -258 0 0 S33
port 68 nsew
rlabel polycont -129 814 -129 814 0 G33
port 69 nsew
rlabel mvpdiffc 0 0 0 0 0 D34
port 70 nsew
rlabel polycont 129 814 129 814 0 G34
port 71 nsew
rlabel mvpdiffc 258 0 258 0 0 S35
port 72 nsew
rlabel polycont 387 814 387 814 0 G35
port 73 nsew
rlabel mvpdiffc 516 0 516 0 0 D36
port 74 nsew
rlabel polycont 645 814 645 814 0 G36
port 75 nsew
rlabel mvpdiffc 774 0 774 0 0 S37
port 76 nsew
rlabel polycont 903 814 903 814 0 G37
port 77 nsew
rlabel mvpdiffc 1032 0 1032 0 0 D38
port 78 nsew
rlabel polycont 1161 814 1161 814 0 G38
port 79 nsew
rlabel mvpdiffc 1290 0 1290 0 0 S39
port 80 nsew
rlabel polycont 1419 814 1419 814 0 G39
port 81 nsew
rlabel mvpdiffc 1548 0 1548 0 0 D40
port 82 nsew
rlabel polycont 1677 814 1677 814 0 G40
port 83 nsew
rlabel mvpdiffc 1806 0 1806 0 0 S41
port 84 nsew
rlabel polycont 1935 814 1935 814 0 G41
port 85 nsew
rlabel mvpdiffc 2064 0 2064 0 0 D42
port 86 nsew
rlabel polycont 2193 814 2193 814 0 G42
port 87 nsew
rlabel mvpdiffc 2322 0 2322 0 0 S43
port 88 nsew
rlabel polycont 2451 814 2451 814 0 G43
port 89 nsew
rlabel mvpdiffc 2580 0 2580 0 0 D44
port 90 nsew
rlabel polycont 2709 814 2709 814 0 G44
port 91 nsew
rlabel mvpdiffc 2838 0 2838 0 0 S45
port 92 nsew
rlabel polycont 2967 814 2967 814 0 G45
port 93 nsew
rlabel mvpdiffc 3096 0 3096 0 0 D46
port 94 nsew
rlabel polycont 3225 814 3225 814 0 G46
port 95 nsew
rlabel mvpdiffc 3354 0 3354 0 0 S47
port 96 nsew
rlabel polycont 3483 814 3483 814 0 G47
port 97 nsew
rlabel mvpdiffc 3612 0 3612 0 0 D48
port 98 nsew
rlabel polycont 3741 814 3741 814 0 G48
port 99 nsew
rlabel mvpdiffc 3870 0 3870 0 0 S49
port 100 nsew
rlabel polycont 3999 814 3999 814 0 G49
port 101 nsew
rlabel mvpdiffc 4128 0 4128 0 0 D50
port 102 nsew
rlabel polycont 4257 814 4257 814 0 G50
port 103 nsew
rlabel mvpdiffc 4386 0 4386 0 0 S51
port 104 nsew
rlabel polycont 4515 814 4515 814 0 G51
port 105 nsew
rlabel mvpdiffc 4644 0 4644 0 0 D52
port 106 nsew
rlabel polycont 4773 814 4773 814 0 G52
port 107 nsew
rlabel mvpdiffc 4902 0 4902 0 0 S53
port 108 nsew
rlabel polycont 5031 814 5031 814 0 G53
port 109 nsew
rlabel mvpdiffc 5160 0 5160 0 0 D54
port 110 nsew
rlabel polycont 5289 814 5289 814 0 G54
port 111 nsew
rlabel mvpdiffc 5418 0 5418 0 0 S55
port 112 nsew
rlabel polycont 5547 814 5547 814 0 G55
port 113 nsew
rlabel mvpdiffc 5676 0 5676 0 0 D56
port 114 nsew
rlabel polycont 5805 814 5805 814 0 G56
port 115 nsew
rlabel mvpdiffc 5934 0 5934 0 0 S57
port 116 nsew
rlabel polycont 6063 814 6063 814 0 G57
port 117 nsew
rlabel mvpdiffc 6192 0 6192 0 0 D58
port 118 nsew
rlabel polycont 6321 814 6321 814 0 G58
port 119 nsew
rlabel mvpdiffc 6450 0 6450 0 0 S59
port 120 nsew
rlabel polycont 6579 814 6579 814 0 G59
port 121 nsew
rlabel mvpdiffc 6708 0 6708 0 0 D60
port 122 nsew
rlabel polycont 6837 814 6837 814 0 G60
port 123 nsew
rlabel mvpdiffc 6966 0 6966 0 0 S61
port 124 nsew
rlabel polycont 7095 814 7095 814 0 G61
port 125 nsew
rlabel mvpdiffc 7224 0 7224 0 0 D62
port 126 nsew
rlabel polycont 7353 814 7353 814 0 G62
port 127 nsew
rlabel mvpdiffc 7482 0 7482 0 0 S63
port 128 nsew
rlabel polycont 7611 814 7611 814 0 G63
port 129 nsew
rlabel mvpdiffc 7740 0 7740 0 0 D64
port 130 nsew
rlabel polycont 7869 814 7869 814 0 G64
port 131 nsew
rlabel mvpdiffc 7998 0 7998 0 0 S65
port 132 nsew
rlabel polycont 8127 814 8127 814 0 G65
port 133 nsew
rlabel mvpdiffc 8256 0 8256 0 0 D66
port 134 nsew
rlabel polycont 8385 814 8385 814 0 G66
port 135 nsew
rlabel mvpdiffc 8514 0 8514 0 0 S67
port 136 nsew
rlabel polycont 8643 814 8643 814 0 G67
port 137 nsew
<< properties >>
string FIXED_BBOX -8906 -952 8906 952
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 7.5 l 1 m 1 nf 68 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 conn_gates 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 doports 1
<< end >>
