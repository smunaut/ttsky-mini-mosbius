magic
tech sky130A
magscale 1 2
timestamp 1756711212
<< metal3 >>
rect 954 27398 1601 27462
rect 1665 27398 1671 27462
rect 0 24310 3680 24610
rect 0 23710 3680 24010
rect 954 22776 1481 22840
rect 1545 22776 1551 22840
rect 0 19688 3680 19988
rect 0 19088 3680 19388
rect 954 18154 1361 18218
rect 1425 18154 1431 18218
rect 0 15066 3680 15366
rect 0 14466 3680 14766
rect 954 13532 1241 13596
rect 1305 13532 1311 13596
rect 0 10444 3680 10744
rect 0 9844 3680 10144
rect 954 8910 1121 8974
rect 1185 8910 1191 8974
rect 0 5822 3680 6122
rect 0 5222 3680 5522
rect 954 4288 1001 4352
rect 1065 4288 1071 4352
rect 0 1200 3680 1500
rect 0 600 3680 900
<< via3 >>
rect 1601 27398 1665 27462
rect 1481 22776 1545 22840
rect 1361 18154 1425 18218
rect 1241 13532 1305 13596
rect 1121 8910 1185 8974
rect 1001 4288 1065 4352
<< metal4 >>
rect 20 27462 260 27550
rect 340 27462 580 27550
rect 660 27462 900 30910
rect 20 22840 260 23110
rect 340 22840 580 23110
rect 660 22840 900 23110
rect 20 18218 260 18488
rect 340 18218 580 18488
rect 660 18218 900 18488
rect 20 13596 260 13866
rect 340 13596 580 13866
rect 660 13596 900 13866
rect 20 8974 260 9244
rect 340 8974 580 9244
rect 660 8974 900 9244
rect 20 4352 260 4622
rect 340 4352 580 4622
rect 660 4352 900 4622
rect 1000 4353 1060 27591
rect 1120 8975 1180 27591
rect 1240 13597 1300 27591
rect 1360 18219 1420 27591
rect 1480 22841 1540 27591
rect 1600 27463 1660 27591
rect 1600 27462 1666 27463
rect 1600 27398 1601 27462
rect 1665 27398 1666 27462
rect 1600 27397 1666 27398
rect 1480 22840 1546 22841
rect 1480 22776 1481 22840
rect 1545 22776 1546 22840
rect 1480 22775 1546 22776
rect 1360 18218 1426 18219
rect 1360 18154 1361 18218
rect 1425 18154 1426 18218
rect 1360 18153 1426 18154
rect 1240 13596 1306 13597
rect 1240 13532 1241 13596
rect 1305 13532 1306 13596
rect 1240 13531 1306 13532
rect 1120 8974 1186 8975
rect 1120 8910 1121 8974
rect 1185 8910 1186 8974
rect 1120 8909 1186 8910
rect 1000 4352 1066 4353
rect 1000 4288 1001 4352
rect 1065 4288 1066 4352
rect 1000 4287 1066 4288
use asw_col_ctrl  asw_col_ctrl_0
timestamp 1756673146
transform 1 0 0 0 1 27598
box -38 -48 3718 3312
use tt_asw_3v3  tt_asw_3v3_0
array 0 0 3680 0 5 4622
timestamp 1756064685
transform 1 0 0 0 1 0
box 0 0 3680 4352
<< end >>
