magic
tech sky130A
magscale 1 2
timestamp 1756676326
<< metal3 >>
rect 1691 19689 1989 19987
rect 1691 10445 1989 10743
rect 1691 1201 1989 1499
<< via3 >>
rect 2291 26763 2589 27161
rect 1691 24311 1989 24609
rect 1691 23711 1989 24009
rect 2891 22141 3189 22539
rect 2291 17519 2589 17917
rect 1691 15067 1989 15365
rect 1691 14467 1989 14765
rect 2891 12897 3189 13295
rect 2291 8275 2589 8673
rect 1691 5823 1989 6121
rect 1691 5223 1989 5521
rect 2891 3653 3189 4051
<< metal4 >>
rect 2290 27161 2590 27162
rect 2290 26763 2291 27161
rect 2589 26763 2590 27161
rect 1690 24609 1990 25462
rect 1690 24311 1691 24609
rect 1989 24311 1990 24609
rect 1690 24310 1990 24311
rect 1690 24009 1990 24010
rect 1690 23711 1691 24009
rect 1989 23711 1990 24009
rect 1690 21240 1990 23711
rect 2290 17917 2590 26763
rect 2290 17519 2291 17917
rect 2589 17519 2590 17917
rect 1690 15365 1990 16218
rect 1690 15067 1691 15365
rect 1989 15067 1990 15365
rect 1690 15066 1990 15067
rect 1690 14765 1990 14766
rect 1690 14467 1691 14765
rect 1989 14467 1990 14765
rect 1690 11996 1990 14467
rect 2290 8673 2590 17519
rect 2290 8275 2291 8673
rect 2589 8275 2590 8673
rect 1690 6121 1990 6974
rect 1690 5823 1691 6121
rect 1989 5823 1990 6121
rect 1690 5822 1990 5823
rect 1690 5521 1990 5522
rect 1690 5223 1691 5521
rect 1989 5223 1990 5521
rect 1690 2752 1990 5223
rect 2290 0 2590 8275
rect 2890 22539 3190 22540
rect 2890 22141 2891 22539
rect 3189 22141 3190 22539
rect 2890 13295 3190 22141
rect 2890 12897 2891 13295
rect 3189 12897 3190 13295
rect 2890 4051 3190 12897
rect 2890 3653 2891 4051
rect 3189 3653 3190 4051
rect 2890 0 3190 3653
use asw_col_base  asw_col_base_0
timestamp 1756676326
transform 1 0 0 0 1 0
box -38 0 3718 30910
<< end >>
