magic
tech sky130A
magscale 1 2
timestamp 1756676326
<< via3 >>
rect 2291 26763 2589 27161
rect 1691 23711 1989 24009
rect 2291 22141 2589 22539
rect 1691 19089 1989 19387
rect 2291 17519 2589 17917
rect 1691 14467 1989 14765
rect 2291 12897 2589 13295
rect 1691 9845 1989 10143
rect 2291 8275 2589 8673
rect 1691 5223 1989 5521
rect 2291 3653 2589 4051
rect 1691 601 1989 899
<< metal4 >>
rect 2290 27161 2590 27162
rect 2290 26763 2291 27161
rect 2589 26763 2590 27161
rect 1690 24009 1990 25462
rect 1690 23711 1691 24009
rect 1989 23711 1990 24009
rect 1690 23710 1990 23711
rect 2290 22539 2590 26763
rect 2290 22141 2291 22539
rect 2589 22141 2590 22539
rect 1690 19387 1990 20840
rect 1690 19089 1691 19387
rect 1989 19089 1990 19387
rect 1690 19088 1990 19089
rect 2290 17917 2590 22141
rect 2290 17519 2291 17917
rect 2589 17519 2590 17917
rect 1690 14765 1990 16218
rect 1690 14467 1691 14765
rect 1989 14467 1990 14765
rect 1690 14466 1990 14467
rect 2290 13295 2590 17519
rect 2290 12897 2291 13295
rect 2589 12897 2590 13295
rect 1690 10143 1990 11596
rect 1690 9845 1691 10143
rect 1989 9845 1990 10143
rect 1690 9844 1990 9845
rect 2290 8673 2590 12897
rect 2290 8275 2291 8673
rect 2589 8275 2590 8673
rect 1690 5521 1990 6974
rect 1690 5223 1691 5521
rect 1989 5223 1990 5521
rect 1690 5222 1990 5223
rect 2290 4051 2590 8275
rect 2290 3653 2291 4051
rect 2589 3653 2590 4051
rect 1690 899 1990 2352
rect 1690 601 1691 899
rect 1989 601 1990 899
rect 1690 600 1990 601
rect 2290 0 2590 3653
use asw_col_base  asw_col_base_0
timestamp 1756676326
transform 1 0 0 0 1 0
box -38 0 3718 30910
<< end >>
